module weight_mat_w2(
	input [31:0] addr,
	output [32*15-1:0] weight
);
	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH = 32;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	32'h3c25ef22,
32'hbdd77885,
32'hbe915f81,
32'h3ead9289,
32'h3e020f09,
32'h3d651423,
32'h3a2a8864,
32'h3f63c5e0,
32'h3ef90cf9,
32'hbdc0a10e,
32'h3f9746f7,
32'h3f27c8f5,
32'hbf5e6fdd,
32'h3faad3be,
32'hbf03b8df,
32'h3e5347b9,
32'hbf3289d9,
32'h3fd5d5a9,
32'h3f56b592,
32'h3eab82f2,
32'h3f099d8c,
32'h3f152e9c,
32'h3f13aa9c,
32'hbee8bec2,
32'h3d25b162,
32'hbf792cc1,
32'hbd38b5ce,
32'h3f199db3,
32'h3f412d51,
32'h3f2b2668,
32'h3e3eb84f,
32'h3f494f4b,
32'h3f10f951,
32'h3e843885,
32'hbd639966,
32'h3e070865,
32'hbcc4cac3,
32'hbd070e39,
32'hbeb8a68f,
32'h3dfd5c9a,
32'hbf550b29,
32'hbe0b99d9,
32'h3f4910d6,
32'h3eb21dac,
32'hbe5fc9c7,
32'h3cdb8e9a,
32'h3deaf2e5,
32'hbe9d019a,
32'h3f18d38d,
32'hbcaa31d4,
32'hbcdcd4ba,
32'hbe1ecf13,
32'hbf2ff789,
32'hbf2a70c1,
32'hbd1a4fb2,
32'hbe8c3838,
32'h3e10d04e,
32'hbe87eb25,
32'hbe3bda14,
32'hbef79252,
32'hbcdfefe5,
32'hbeee0e2b,
32'h3f49d8f1,
32'h3f029a1d,
32'h3d1e6dee,
32'h3dd500f3,
32'h3d81c372,
32'h3e1825ab,
32'hbee6b244,
32'hbeace7a1,
32'h3f1d5cea,
32'h3f00b63e,
32'hbafbdff1,
32'h3e94a637,
32'hbe079915,
32'h3c1255d9,
32'hbddf35ac,
32'hbee86b57,
32'h3eafcd21,
32'hbca96208,
32'hbf9bdb48,
32'h3ded68aa,
32'h3ee90c3f,
32'h3f1e778c,
32'hbdbff698,
32'h3f164fd4,
32'hbc1a6075,
32'hbf2a2f1c,
32'h3f5a75c4,
32'hbe95cbdd,
32'h3d80c3a4,
32'h3dc384aa,
32'h3ec2f15a,
32'hbeffade7,
32'hbd22ab21,
32'h3c877be7,
32'h3d30481c,
32'hbf11f5ed,
32'hbe6399a1,
32'h3dbaa969,
32'hbe95626d,
32'hbe98e75d,
32'h3eae4d90,
32'hbddbdf0a,
32'h3f232dfa,
32'h3d28a5ce,
32'h3d8bb51e,
32'h3f23f6bd,
32'h3e91ba34,
32'hbdcd577b,
32'hbd26a415,
32'h3e673d3c,
32'hbef7371d,
32'h3ec992ce,
32'h3d62a246,
32'hbe025cfc,
32'hbef5eccf,
32'hbe4af8ed,
32'hbea9718c,
32'h3f4242ca,
32'h3ea83225,
32'h3f8b37c9,
32'h3e9374cd,
32'h3e28e0ab,
32'h3bbb0dd0,
32'h3e2014f9,
32'h3d11d38e,
32'h3ecb03f5,
32'h3dd8280f,
32'h3f244b61,
32'hbfc06298,
32'hbf36f1ec,
32'h3f994fb8,
32'h3e7e5008,
32'h3e8b7ae2,
32'h3d797de3,
32'h3eb4ca4f,
32'hbf9b129f,
32'h3dcaca48,
32'h3e09171b,
32'h3d2fb713,
32'hbdc165a1,
32'h3f579007,
32'hbf3ba61c,
32'h3d009fa4,
32'h3f5e9585,
32'h3eb8c97a,
32'hbe169c2b,
32'h3f9b5fce,
32'hbf5da521,
32'hbd7daa61,
32'h3e69fc85,
32'h3f10508c,
32'h3e430603,
32'hbd3c8730,
32'h3e135366,
32'hbe4077c8,
32'hbee30e12,
32'h3e7941cc,
32'hbf0b7e99,
32'h3d8de9b2,
32'h3e63caa3,
32'h3d166b4b,
32'hbea7f2cc,
32'h3d01602d,
32'h3ed4d069,
32'h3e44463d,
32'hbcc78930,
32'h3c03f1d2,
32'hbd2aa3d4,
32'h3e64125e,
32'h3e636228,
32'h3d8edb59,
32'hbd861b0b,
32'h3e2bb2e2,
32'h3e88274f,
32'hbe3f34ba,
32'hbeac06c3,
32'h3ca1922d,
32'h3b6e7ad0,
32'hbc91c987,
32'h3e1d6e82,
32'hbf417e98,
32'h3e2775d4,
32'hbf001202,
32'hbde4abfb,
32'hbe4dfd38,
32'hbead31cb,
32'h3e87fb4b,
32'hba9d66d9,
32'hbccf5d29,
32'hbe48a528,
32'h3ed99a76,
32'h3e4787c6,
32'hbea0ca73,
32'h3e831f92,
32'h3f86334f,
32'hbe8165ec,
32'hbf6f23b5,
32'hbeb3ec64,
32'h3dd70927,
32'hbdc1231d,
32'h3e6dcaaf,
32'hbd867aa2,
32'h3f02d2c0,
32'hbe215605,
32'hbf16d7c9,
32'h3fbd9fec,
32'h3f0186da,
32'hbe05847a,
32'h3e355ffc,
32'h3f300c55,
32'h3e13b757,
32'hbefd513c,
32'hbd50f309,
32'h3e070be5,
32'h3d029504,
32'h3eb91594,
32'hbd5fcbc2,
32'h3eb50b5a,
32'hbe843978,
32'hbe9bb95d,
32'h3f23e27b,
32'h3f446265,
32'h3e57327a,
32'h3bb27b9d,
32'hbe76b85e,
32'hbeb78506,
32'hbe02f594,
32'h3d01fbb6,
32'hbbc88f26,
32'hbd3f8d7f,
32'h3e356461,
32'hbf4278ae,
32'h3d299c51,
32'hbec37052,
32'hbd1345c2,
32'hbd5a1347,
32'hbe4fc568,
32'hbce9b764,
32'h3e7aed24,
32'h3f750661,
32'hbf556f4a,
32'hbeffe5df,
32'hbe05fdb2,
32'hbdd41f8d,
32'hbd4904f8,
32'h3e69300f,
32'hbf6c41fe,
32'h3f046a34,
32'h3eb415fb,
32'hbe0bf9d4,
32'h3f07a9bc,
32'h3f200d24,
32'hbe4b4070,
32'hbd1f8815,
32'h3d0ed2b8,
32'hbfb36087,
32'hbf8b5a69,
32'hbe863179,
32'h3e263dff,
32'hbe9f186e,
32'hbf2abf2b,
32'hbe990511,
32'hbe9e313f,
32'h3e292a35,
32'h3f5d131d,
32'h3ec72f93,
32'h3f1ce7e5,
32'hbf0816e0,
32'hbd1781ae,
32'hbeec59ec,
32'h3f28f844,
32'h3eb26f74,
32'h3dabd011,
32'h3d4089fe,
32'h3da31c3e,
32'hbe460596,
32'hbea36724,
32'hbe96f2ff,
32'h3ecfd208,
32'h3e4f47ea,
32'hbe4397c0,
32'hbda044e6,
32'hbecb1a1b,
32'hbd91e7b0,
32'hbee7f5ca,
32'hbe1f8214,
32'hbef5ac95,
32'h3cb6bb99,
32'h3e373de4,
32'hbc4152d1,
32'hbe8cdcb2,
32'h3ec15de3,
32'hbed2e6c1,
32'h3f12597a,
32'h3f2f246c,
32'h3e1815d6,
32'h3e8e3889,
32'h3e778578,
32'hbd757cfd,
32'hbd84def5,
32'hbf502920,
32'hbf2dbb38,
32'hbe183986,
32'h3e273252,
32'hbde55ad8,
32'hbf50fe47,
32'hbeea3c34,
32'hbeed5cf9,
32'h3ecb1310,
32'h3f1fe341,
32'h3ef8ce9e,
32'h3e6a844d,
32'hbf14be5b,
32'h3bcc4b49,
32'hbead114e,
32'hbf240cfd,
32'hbe9a31a0,
32'hbb5de868,
32'h3ac10e3d,
32'h3cac33bf,
32'hbeeba4f2,
32'hbd521bc8,
32'hbc95e25c,
32'hbf09c0e0,
32'hbe427766,
32'hbf4c75da,
32'hbf2d6905,
32'hbe918bfc,
32'hbeeaa14c,
32'hbf227b57,
32'h3f181be6,
32'h3e9875bf,
32'hbf846ee9,
32'hbf242b96,
32'hbe95567f,
32'hbfca8a10,
32'h3ec1a6fc,
32'hbf8c54c9,
32'hbf5b7b38,
32'hbed4b519,
32'h3f396e5c,
32'hbf448fce,
32'hbf67baa7,
32'hbc5cdf91,
32'hbd59a359,
32'hbdb1f1a4,
32'hbdcf8c51,
32'hbd32c7a4,
32'hbca8ad50,
32'hbbeb2660,
32'hbe7df495,
32'hbf03a693,
32'hbdad9564,
32'hbe90181d,
32'hbe6fca06,
32'h3d7d90f7,
32'hbedf886c,
32'hbf13f17f,
32'h3dc4ded1,
32'h3e6ec3a1,
32'h3f135a42,
32'h3e0e63f5,
32'hbd170a0a,
32'h3d056092,
32'h3e00b9d3,
32'hbea19ece,
32'h3dc2f084,
32'h3db9670d,
32'hbf42d175,
32'hbe2bf50b,
32'h3e8a1fd4,
32'hbd2e4173,
32'h3f428526,
32'h3e2e0024,
32'hbed58f47,
32'h3f7a734c,
32'h3f31f942,
32'h3e245ee8,
32'h3ed0f118,
32'h3eb6c98f,
32'h3ee2cdb9,
32'hbef61837,
32'hbdd6eb34,
32'hbf15a645,
32'h3d78c4b0,
32'h3ec5a214,
32'h3ecb6bb7,
32'h3e963b8b,
32'hbaaf65b4,
32'hbdc05069,
32'hbebef5b9,
32'hbe68db09,
32'hbb81871b,
32'hbd55d4a4,
32'h3a4a42a9,
32'hbe3fb262,
32'h3e81f9ec,
32'h3cbe3ec1,
32'hbe1ea538,
32'hbf10371b,
32'hbe3e6ae4,
32'hbf01e152,
32'h3d8ecbb2,
32'h3a2c2ee4,
32'hbdaba94a,
32'hbe99adde,
32'hbe8280dd,
32'hbdc33526,
32'hbf998c0b,
32'h3e64afce,
32'hbf9f2282,
32'h3f91aa3b,
32'hbde78fce,
32'h3e5ad414,
32'hbfd788d8,
32'hbe90675c,
32'h3c3ca1e7,
32'h3d3a9628,
32'h3e5acb4e,
32'h3f313668,
32'hbe59ca3f,
32'hbe0ccf34,
32'hbf413dea,
32'hbd417091,
32'hbc910af4,
32'h3e901ec1,
32'hbedce184,
32'h3f36d266,
32'h3e886198,
32'hbf2f7999,
32'h3f9658d8,
32'h3f19f43f,
32'h3ef233b7,
32'hbd058e57,
32'h3c8ab14d,
32'hbe83cc8e,
32'hbf0985bf,
32'hbdd60cfa,
32'h3cdea670,
32'hbe05a1b8,
32'hbe4a4a40,
32'hbe588fee,
32'hbd9349ce,
32'hbf4aff83,
32'h3e3c8059,
32'hbf02d1f9,
32'hbeb7417b,
32'hbe8af785
};
	assign weight = {ROM[addr],ROM[addr+1],ROM[addr+2],ROM[addr+3],ROM[addr+4],ROM[addr+5],
						ROM[addr+6],ROM[addr+7],ROM[addr+8],ROM[addr+9],ROM[addr+10],ROM[addr+11],
						ROM[addr+12],ROM[addr+13],ROM[addr+14]};

endmodule 