module weight_mat_w1(
	input [31:0] addr,
	output [32*30-1:0] weight
);
	parameter ADDR_WIDTH = 15;
   parameter DATA_WIDTH = 32;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	32'hbcd6c54c,
32'h3d821706,
32'h3d317bf2,
32'hbcdd0db5,
32'hbd88d9f1,
32'hbc463af5,
32'hbd1e508c,
32'hbc22ac22,
32'hbd468956,
32'hbd7d7352,
32'hbc7f0974,
32'h3d631565,
32'h3d97a41a,
32'hbd4e33cc,
32'hbd833006,
32'h3ce94a1d,
32'hbd0180de,
32'hbd3b8610,
32'hbd19378e,
32'h3c7c5fc3,
32'h3ca58c5a,
32'hbd1f4833,
32'h3d03bf1f,
32'hbb7d6ea0,
32'h3c8cd1b1,
32'hbd9d7a36,
32'h3ce32247,
32'hbd85476b,
32'hbc137ea0,
32'hbc2c2f07,
32'h3b585e25,
32'h3cd1ec07,
32'hbc0f8ff9,
32'h3d53a11e,
32'h3d1590ed,
32'h3d541b34,
32'hbd9aeec4,
32'hbd9a893a,
32'hbade29c0,
32'hbd51be02,
32'h3bf052e7,
32'hbdb42158,
32'h3d9bfecf,
32'h3cff9868,
32'h3dba8036,
32'hbca06f44,
32'h3dc20bb9,
32'h3ca1f580,
32'hbd6a5644,
32'h3bb8cc8d,
32'hbd9825f1,
32'hbcfd9974,
32'hbca783a8,
32'hbd2d360d,
32'h3d84a97b,
32'hbcd2a216,
32'h3cbf45da,
32'hbce36a1d,
32'hbd1b94ac,
32'hbcd4b4cc,
32'h3dbecf72,
32'hbccafb28,
32'hbd30fab0,
32'h3c85a312,
32'h3d75a0d4,
32'h3cff1df7,
32'hbd8f849b,
32'hbca140ca,
32'h3c8c5eaf,
32'hbd97abc4,
32'hbce673a0,
32'h3d4af725,
32'h3c85dbf3,
32'h3db529f7,
32'h3d9a2030,
32'hbce8f1e5,
32'h3d2c11c7,
32'hbc27f4bd,
32'hbc9a0244,
32'h3de049ed,
32'hbc3ca6cf,
32'hbd98ac79,
32'h3d1a4ae2,
32'hbce8c7e2,
32'h3c71e4f4,
32'h3d7417a1,
32'hbd583ade,
32'h3d77f2a6,
32'h3ca7ce9a,
32'h3d09c21d,
32'h3d65d628,
32'hbc9c954f,
32'h3d17f2b1,
32'hbbc579f6,
32'hbd396cdd,
32'h3d32fddd,
32'hbdd07080,
32'h3db99cb0,
32'h3c824155,
32'hbd90c993,
32'h3d33b07a,
32'hbdbbf1f2,
32'hbc2e9691,
32'hbd7b5dcb,
32'hbd0da511,
32'h3ccf553a,
32'hbd7c241b,
32'hbd837dac,
32'h3db9c066,
32'hbd1fba45,
32'h3ca4d1cc,
32'hbc816f00,
32'hbc21cf4f,
32'h3d64ba0b,
32'h3d177d50,
32'hbdad3e96,
32'h3d1e3918,
32'h3d617b6d,
32'h3d7fda78,
32'h3d608f17,
32'hbc9c714f,
32'h3d644a7e,
32'h3d7f2cda,
32'h3cc35d65,
32'h3c99da2a,
32'hbd19717c,
32'h3c8431ad,
32'h3ae55f51,
32'hbd98d8dc,
32'hbc54207a,
32'hbcb5cf50,
32'hbdac8193,
32'hbd9486e1,
32'hbd09f692,
32'hbc9d64db,
32'h3b98c91c,
32'hbd412c64,
32'h3cbde416,
32'h3d06e87c,
32'h3dbe1b49,
32'h3b959ec3,
32'h3c7b535d,
32'h3d2760b9,
32'h3d1211a9,
32'hbbe2a23f,
32'hbdb989b2,
32'hbd27b3bb,
32'h3cf5f2eb,
32'hbd1b2545,
32'h3d5f9af2,
32'hbd881115,
32'h3cbd435b,
32'hbcbe5691,
32'h3c0023cb,
32'h3d71ab48,
32'h3d6ef53a,
32'h3b208619,
32'hbd7530b0,
32'hbcca41f1,
32'hbd92e122,
32'hbd8d0993,
32'hbd2f7da9,
32'h3d8e1043,
32'hbd66732e,
32'h3d493955,
32'hbd3862dd,
32'hbd104c9a,
32'h3cc7fcaf,
32'h3c5cef08,
32'h3c3d1226,
32'h3c80b1f6,
32'hbdcb99b4,
32'hbc895476,
32'hbd51a559,
32'h3cf8ef65,
32'h3c6e9847,
32'h3c5c3bc3,
32'hbb8b8965,
32'hbc65e19c,
32'hbd9aff00,
32'hbd770b62,
32'h3bf26b73,
32'hbd429e58,
32'hbb8bba3e,
32'h3bdbaa89,
32'hbcc4e5ea,
32'h3d2f3c1c,
32'hbb58293f,
32'hbd98cc97,
32'h3b83ab27,
32'h3b95b48b,
32'hbd33a073,
32'hbd88aa27,
32'hbacc6118,
32'hbbd3cce1,
32'h3c8239bd,
32'h3cd2057c,
32'hbcb18eb4,
32'hbb3b0dd9,
32'h3dc6efe9,
32'h3d282b97,
32'h3d66f3e9,
32'hbc3b9310,
32'hbd245f88,
32'h3d530da3,
32'hbcbdb363,
32'h3d973bb8,
32'hbcf51341,
32'h3b2d6071,
32'hbda83505,
32'hbd70891b,
32'h3db0b015,
32'h3d25dff9,
32'h3dce6ee0,
32'h3c98a258,
32'hbc23ccd5,
32'hba1a1cc8,
32'hbd186e5a,
32'hbcb07135,
32'h3d839e08,
32'h3d770136,
32'h3c2a8a8a,
32'hbda469b9,
32'h3d1187f6,
32'h3d9e5147,
32'hbd6882f1,
32'h3d2c1600,
32'hbdb3fc02,
32'h3d33e1e1,
32'h3c8150a2,
32'hbd8843b1,
32'h3d3890c5,
32'h3d3d9cce,
32'h3d52432e,
32'hbc63c99c,
32'hbbc97a31,
32'h3d03bb6a,
32'h3cfda2d2,
32'hbc5a8786,
32'h3d71d034,
32'h3d00694e,
32'h3cb0c885,
32'hbd9c3154,
32'h3d89a0d3,
32'h3d273d72,
32'h3c14fd4c,
32'h3d5f8900,
32'hbc21c7b3,
32'hbc88f40e,
32'h3cb63773,
32'h3d0b4116,
32'h3d44d4e5,
32'h3d6a634e,
32'hbd03c020,
32'hbdd96144,
32'h3d9223ac,
32'h3db418d6,
32'h3d5ae39e,
32'hbcda0c6a,
32'hbc4c07b7,
32'hbcab3614,
32'h3c14c439,
32'h3c8ffcc3,
32'hbd38e3ce,
32'hbbebb8f3,
32'hbcb6ed9e,
32'hbba877e5,
32'h3dad81b3,
32'h3d9e5acb,
32'h3d4c5861,
32'h3c8c6fda,
32'h3d890d95,
32'hbbb9a8cd,
32'hbd02a3ab,
32'hbd010dbf,
32'h3cae5a34,
32'hbcc23ab0,
32'h3c2e9b2b,
32'h3d929446,
32'h3da2dd81,
32'h3d31a91f,
32'h3d14b720,
32'h3d2eeb78,
32'hbd8c95d6,
32'h3c97acfe,
32'h3d89a9d7,
32'hbc62db39,
32'h3d577e93,
32'hbcb3d837,
32'hb93b3124,
32'hbd102f28,
32'h3cce54f4,
32'h3de9a9ac,
32'h3d0ef741,
32'hbce2e454,
32'h3d5e83ef,
32'h3be35399,
32'hbc62cbed,
32'h3ac6f5d0,
32'hbdace555,
32'hbc707538,
32'h3c8684c8,
32'h3d486886,
32'hbd3f6594,
32'h3d50979c,
32'h3d12db26,
32'hbd96e718,
32'h3d37de34,
32'h3d1b2a3c,
32'hbd3756b6,
32'hbcade987,
32'h3d575b60,
32'hbdaf59d6,
32'h3d6e5c3f,
32'h3dcceee9,
32'h3cf4c268,
32'hbd4fe6fe,
32'hbd84df8f,
32'h3cb9d9f3,
32'hbd2b34a4,
32'hbd4927a7,
32'hbc9d04c9,
32'h3c9a1579,
32'hbb39d9a7,
32'h3b88e2d9,
32'h3c93d566,
32'hbc9ed878,
32'h3d074571,
32'hbdb259c4,
32'hbd0856fd,
32'hbbea0b68,
32'hbc6c65f8,
32'hbd228510,
32'h3c14e635,
32'h3d4ebcf0,
32'hbc0ddf21,
32'hbcf5f551,
32'h3c1d93f7,
32'h3db56678,
32'hbbf919ef,
32'hbdda5bcb,
32'h3d7ec61d,
32'hbd089994,
32'hbda7ecea,
32'hbcb00954,
32'hbc8abd6d,
32'hbd8b2c3a,
32'h3d1c321c,
32'h3d02ac2a,
32'h3d936a8d,
32'h3c962a06,
32'h3d139ddb,
32'hbcc3ba55,
32'hbd0f4e59,
32'hbd2d1c6f,
32'hbdaec6a1,
32'hbbf6dfe9,
32'hbc056b16,
32'h3dd99a26,
32'hbd8e9e05,
32'hbdb57a76,
32'hbb1d0f3c,
32'h3c94355b,
32'hbdab8c4f,
32'hbb5d856b,
32'h3d468168,
32'h3d8bff51,
32'h3d29377e,
32'h3a6b1938,
32'h3d8a48c5,
32'hbcbed7fe,
32'h3acad110,
32'hbd67b716,
32'h3e275058,
32'h3cfb2f37,
32'hbcef304e,
32'h3cbae6e1,
32'hbd1bf540,
32'h3da7b86a,
32'hbd6bff55,
32'h3d86025a,
32'hbdfe10d5,
32'h3cc00afd,
32'hbe1a0316,
32'h3d7eaec0,
32'h3cbb14d9,
32'h3e1b11ce,
32'h3ccc0fa8,
32'h3b418c60,
32'hbd8b9ea8,
32'h3db2d916,
32'hbd3b25ed,
32'h3ca7c815,
32'h3c6defde,
32'hbda92315,
32'h3c706f6b,
32'h3d86c094,
32'h3a0ef35c,
32'h3d6aa13a,
32'hbd43e053,
32'hbc03be84,
32'h3db6a4a3,
32'h3bba85fe,
32'h3dfaa419,
32'h3e1a8ea5,
32'hbe51fbc8,
32'hbd615cd9,
32'h3c750650,
32'h3cdb2c20,
32'h3ceb540c,
32'h3ca8d5ae,
32'hbe291810,
32'h3d2dae13,
32'hbe856aca,
32'h3e68cd9b,
32'h3d04bce8,
32'h3e3b32c1,
32'hbda143f6,
32'h3e3bb1ef,
32'hbdcdef4a,
32'hbcd019ca,
32'hbcd6382f,
32'hbc11e363,
32'h3c049ba6,
32'hbdb00c1e,
32'h3cfc8880,
32'hbd831f76,
32'h3d38f79e,
32'h3e21a882,
32'h3d4bbb18,
32'h3d223879,
32'h3de13f23,
32'h39d5cc62,
32'h3e153fce,
32'h3e6621b6,
32'hbe147444,
32'h3c959078,
32'hbd554d43,
32'hbd288d1e,
32'hbc6d44eb,
32'hbdcb874b,
32'hbe1ed1c5,
32'hbd926626,
32'hbe6cfb2a,
32'h3e5d2403,
32'hbdb04840,
32'h3e33ca15,
32'hbd0be0d4,
32'h3ce0e0a2,
32'hbc914540,
32'h3d530dad,
32'hbda1e32c,
32'hbc11ba56,
32'h3cda6cf6,
32'h3d00e169,
32'h3d091f4f,
32'hbd82c82e,
32'h3d2f4804,
32'h3dead0f4,
32'hbd5affbb,
32'hbc8ef8b4,
32'h3d7b212c,
32'hbcbe5ba8,
32'h3de76e04,
32'h3c288896,
32'hbd55e055,
32'h3d7af44e,
32'h3c875ac5,
32'h3d9e8a52,
32'h3de0c319,
32'hbcc30055,
32'hbda7db04,
32'h3d845f24,
32'hbe2bce63,
32'h3b821e70,
32'h3cba27e9,
32'h3d68802d,
32'h3d9c27cf,
32'h3bd91897,
32'hbd20a49e,
32'h3c7966eb,
32'hbd45ac45,
32'hbd97aaf3,
32'hbdce106b,
32'h3c827e57,
32'hbd968324,
32'h3c552137,
32'h3d727959,
32'h3c3f4383,
32'hbd96c57f,
32'hbceceffe,
32'h3db7852e,
32'hbc9e84df,
32'h3dcda38c,
32'h3d460b35,
32'h3d9c867f,
32'h3dde16bc,
32'h3c6a4055,
32'h3d59425c,
32'h3d32fedd,
32'h3ce63ec0,
32'h3d013239,
32'h3d6dfda4,
32'h3d138cec,
32'h3cfb30e9,
32'hbd89a3dd,
32'h3bfafeaf,
32'h3d6ddde3,
32'hbcd5f923,
32'hbc83dbdd,
32'h3cdeedae,
32'hbd8b4fb5,
32'hbca65c99,
32'h3c6936cb,
32'hbbfce99d,
32'h3c7b3de1,
32'hbd5592b2,
32'hbbbbda4c,
32'hbcbbcb4e,
32'h3cc9ed9b,
32'hbc14b3c7,
32'h3cdb1e96,
32'hbbae7159,
32'h3d43107f,
32'h3de8b3e4,
32'h3c0c0e96,
32'h3cafeaf5,
32'hbdbd1566,
32'h3b2342b4,
32'hbdbeb34a,
32'hbd62e92d,
32'hbcaf1658,
32'hbcb8e371,
32'hbd1fece5,
32'hbd3b75b1,
32'h3cfa04c7,
32'hbd156310,
32'hbcbda790,
32'hbd26e8d6,
32'hbcbe0c73,
32'hbcfa516a,
32'hbca40db2,
32'hbcc5f040,
32'h3d4efeb2,
32'hbcf49742,
32'h3b15c376,
32'hbd8def06,
32'h3c3fb94f,
32'hbd8d3125,
32'hbb5aea65,
32'h3d5f1452,
32'hbdbb64e5,
32'hbd30edcf,
32'hbd62748f,
32'h3d368525,
32'h3d00bfa2,
32'h3d5f6ad2,
32'hbc27a076,
32'h3d8e39d1,
32'hbc5b9873,
32'h3cb60d36,
32'hbdc016ad,
32'hbb86f6d0,
32'hbd0472d2,
32'h3c19c924,
32'hbd497af8,
32'hbd4e34aa,
32'hbd71b6cf,
32'hbb6cadd8,
32'hbc503baa,
32'h3bd4d34a,
32'hbb25f1c1,
32'h3c260b04,
32'h3d9a26dc,
32'h3c8a6684,
32'hbd86d099,
32'hbd99153e,
32'hbd565daf,
32'hbd671f81,
32'h3d647e45,
32'hbd44afcf,
32'hbd11d7f6,
32'hbb271759,
32'hbd917920,
32'hbc9bc2ec,
32'hbbfdd64f,
32'h3c8f2831,
32'h3dba300d,
32'h3d9d49ca,
32'h3d666700,
32'hbd252948,
32'hbdacc1fe,
32'h3d323ca7,
32'hbbb9b38e,
32'hbd27649a,
32'h3d8f757b,
32'hbd46e2d0,
32'h3dad2adf,
32'hbd1a0142,
32'hbdb4d6da,
32'h3d115267,
32'h3c65c81d,
32'h3c8cab5f,
32'hbd4ff9af,
32'h3dcc21c9,
32'h3b5c0190,
32'hbd21a54a,
32'h3d4f224a,
32'hbd013ee2,
32'hbcda853f,
32'hbd21d42b,
32'hba485720,
32'hbdd95682,
32'h3d32907b,
32'hbd984f67,
32'h3ceafd62,
32'hbc9fc67b,
32'h3be294f1,
32'h3d268a38,
32'hbd78280a,
32'h3d19cc32,
32'h3c4fec95,
32'h3d1127bf,
32'hbd5e4d54,
32'hbdbcabc6,
32'h3c4bbab8,
32'h3dce0031,
32'h3a85f07e,
32'hbc8d4bcd,
32'h3d0a1531,
32'hbb87b492,
32'h3d96b0ad,
32'h3c64b66f,
32'h3d4a52cb,
32'h3caf26a7,
32'hbdd891d6,
32'hbccb777b,
32'h3cd826f7,
32'hbd85dd54,
32'h3dc30776,
32'hbd29cbb4,
32'hbc80b6f7,
32'hbd9816b1,
32'h3d86303d,
32'hbd31cafc,
32'h3c0f8313,
32'h3bf56e8f,
32'h3ceb6a68,
32'h3c54eb65,
32'h3d69b9b3,
32'h3d643108,
32'h3ce5b55f,
32'h3d4e51de,
32'hbcbda9f5,
32'hbcb4d4bc,
32'h3c4da178,
32'hbd0fb7c2,
32'h3d4d0705,
32'hbd699243,
32'h3d0d2869,
32'hbd344717,
32'hbcea6eec,
32'h3bdb574c,
32'hbc64863d,
32'hbb4c55b7,
32'hbcab6873,
32'h3cb0883f,
32'h3c00a28f,
32'h3cff8dcc,
32'hbbeb7878,
32'h3cb51746,
32'hbccd4070,
32'hbd7a6853,
32'hbdd31aea,
32'hbbef770d,
32'h3d4d8b51,
32'h3b8c7472,
32'hbdc01c6e,
32'hbd36e64c,
32'h3d2288a7,
32'h3d353345,
32'h3dc40d7d,
32'h3c24918e,
32'hbd4ba5b4,
32'h3dde09b7,
32'hbc5bc926,
32'hbcebe371,
32'hbc861b81,
32'hbd9923df,
32'h3d9e2619,
32'hbc8e8fce,
32'h3a6c0e6d,
32'h3d263a58,
32'hbad03cff,
32'h3c888f49,
32'hbd02bbbb,
32'hbd6f8e24,
32'hbd3ba317,
32'h3d9170ad,
32'h3c962db7,
32'hba9412df,
32'h3c8b80a7,
32'h3c85faba,
32'h3d7bc6cc,
32'hbd25a3e1,
32'h3d203f06,
32'hbbd492a9,
32'h3d7ddeb9,
32'h3da597d6,
32'h3d3ca7cb,
32'hbda535e9,
32'h3d3f9dee,
32'hbcb142eb,
32'h3dc21533,
32'h3d114f7d,
32'hbd051384,
32'h3cae3a89,
32'h3d7f2b91,
32'hbca5449f,
32'h3cafce81,
32'hbcf21d4e,
32'h3dcc28bd,
32'h3db6bfa6,
32'h3bf4349c,
32'h3d002ad6,
32'hbc5db306,
32'hbab3d63f,
32'hbc699b55,
32'h3d237eaf,
32'hbcf2ca42,
32'h3d46420d,
32'hbd668a30,
32'hbd1ff62a,
32'hbb6f0d0e,
32'h3d39561c,
32'hbd170854,
32'hbd500703,
32'h3dcd6bec,
32'h3c7dfdba,
32'hbcb6ffc7,
32'hbc34d51b,
32'hbc0025e4,
32'hbc544719,
32'hbd9b3686,
32'h3c9d10e8,
32'h3abd9569,
32'hbc05fd0e,
32'hbc943aef,
32'h3c319a7c,
32'h3ccb560e,
32'h3ca014d8,
32'h3d81a7f1,
32'h3c1b04bc,
32'hbc6bc8a4,
32'hbd23566f,
32'hbdd26dea,
32'hbc0f940b,
32'hbc775925,
32'h3da99615,
32'hbd3174f7,
32'h3d75a584,
32'hbd86926c,
32'h3c7fa14d,
32'hbd186b3f,
32'h3d1d0ed0,
32'h3d0b4619,
32'h3d20e89e,
32'hbd994897,
32'hbc718456,
32'h3c34ca03,
32'h3cc68697,
32'hbd02f393,
32'hbca97a02,
32'hbd9a527a,
32'h3d0f4d54,
32'h3dd803c5,
32'hbd947719,
32'hbd52fe16,
32'hbdc9dd5a,
32'h3cb9a14b,
32'h3daabc99,
32'h3cd0e75a,
32'hbc508d75,
32'hbc277def,
32'h3bf47459,
32'hbb9fce99,
32'hbd61ddba,
32'h3d2eefac,
32'hbc18d627,
32'h3c89a2dd,
32'h3cb1bc89,
32'h3cdf828e,
32'h3d6a5048,
32'h3d215419,
32'h3da5d48e,
32'hbc796f35,
32'h3dbd28bd,
32'h3bd804b8,
32'hbb755df9,
32'h3d8ca12b,
32'hba924daa,
32'hbd22b249,
32'hbd7594fd,
32'hbc394124,
32'hbd2ed32a,
32'h3d7f0063,
32'hbd170ad0,
32'h3d77bdc2,
32'hbdaf259a,
32'hbdd99341,
32'hbd23b33f,
32'h3d3e20e1,
32'hbd816ada,
32'h3ab67f2c,
32'h3d3f5df8,
32'h3c439a1d,
32'h3cbd899d,
32'hbcb04b72,
32'hbcad2dd0,
32'hbd3fd60c,
32'hbd03f957,
32'h3d8083c4,
32'hbd1023bf,
32'h3d93c925,
32'h3d3f077e,
32'hbcceb515,
32'hbdac33f4,
32'hbd13d20f,
32'hbc8ee2f0,
32'hbca33573,
32'hbdbefa28,
32'hbd7267fc,
32'hbd171ffb,
32'hbcd21c8a,
32'hbd57f0c3,
32'hbd54e136,
32'hbd44e526,
32'hbb7418e6,
32'hbddc9871,
32'hbd07c8f1,
32'h3d217482,
32'h3d5cb472,
32'hbc34fb82,
32'h3d516051,
32'h3d61c33b,
32'h3dbe4258,
32'h3d8533a8,
32'hbdb237fb,
32'hb9637ddc,
32'hbd7239a0,
32'h3d6174d3,
32'h3d3bcd6d,
32'hbcbea41d,
32'hbd5fed8c,
32'hbd2b4c5f,
32'hbcf76d57,
32'h3b33caec,
32'h3c0cb334,
32'h3d205361,
32'hbcbec5bb,
32'h3cb70a3c,
32'h3cdb1e2b,
32'h3ddb88d9,
32'h3d65091c,
32'h3dc478e1,
32'h3d29382b,
32'hbd0815fc,
32'h3c6d5bf8,
32'h3daf695d,
32'hbc825300,
32'h3da4ce29,
32'hbcc71f3e,
32'hbd2341fb,
32'h39940659,
32'hbc7c05b5,
32'hbc59c42c,
32'hbc1b6b7f,
32'h3d877476,
32'h3db1eb40,
32'hbdb6696d,
32'h3d25f87a,
32'h3da68bc7,
32'h3d75a891,
32'h3cd8e1d4,
32'h3d201736,
32'h3d218b3a,
32'hbcdbc661,
32'hbdbf0cc1,
32'hbcf81041,
32'hbd65059c,
32'h3d1998bd,
32'h3d35f5f0,
32'h3dc4aeca,
32'h3d11384b,
32'hbd377a0c,
32'hbbcf3e0c,
32'hbcbcca83,
32'h3d401625,
32'hbd234366,
32'h3c8d24de,
32'h3ca20145,
32'hbcae0ac3,
32'h3d3085a4,
32'hbca36fc1,
32'hbd8a80b9,
32'h3d98e0aa,
32'hbc8b5e83,
32'h3c0d1fb3,
32'hbb98a05c,
32'h3c8fc03b,
32'h3d23f38a,
32'hbd2399a8,
32'h3d317e56,
32'hbcef6888,
32'h3c6a5fef,
32'hbc313f25,
32'hbcd9059e,
32'h3c676b90,
32'h3d3a58f7,
32'hbcb9323a,
32'h3b3d2add,
32'hbdc77c16,
32'hbcb2128d,
32'h3a690bb3,
32'h3d167396,
32'h3cf3b862,
32'h3da3e147,
32'h3d3038e8,
32'h3c1f4f61,
32'h3de7976b,
32'h3c8894f0,
32'hbb60e470,
32'h3dacf5f2,
32'h3cdae3c3,
32'h3c88277f,
32'h3d1c006c,
32'hbdb68ae6,
32'h3d45d698,
32'hbd50e14e,
32'hbd5c3961,
32'hbb2ff790,
32'h3d273901,
32'h3c73552f,
32'hbde47016,
32'hbd8541a1,
32'hbd3410c0,
32'h3c8f6340,
32'h3dae81b0,
32'h3c7d68a3,
32'hbcac29ea,
32'hbcc0f763,
32'h3c9797df,
32'hbdcdeb50,
32'hbb88ace7,
32'h3c9a533d,
32'hbbcd98ba,
32'h3d77415d,
32'h3d118941,
32'h3d45c952,
32'h3dcb3289,
32'hbd2a8866,
32'h3d4869d7,
32'hbdb3168c,
32'h3c89ea44,
32'hbde42e5b,
32'h3da6d07d,
32'hbd79b8e6,
32'hbcc1c891,
32'hbcdc17c1,
32'h3d539edf,
32'hbbc2399d,
32'hbd3512c2,
32'h3cda5726,
32'h3c8842a6,
32'h3d2b53df,
32'hbcda2613,
32'hbb016ab4,
32'hbd8a0ddd,
32'hbcc7e027,
32'hbd07dca9,
32'hbc559915,
32'h3d4bcb99,
32'hbd268b06,
32'h3d4c5392,
32'h3ddd3ddf,
32'h3ad7d229,
32'hbcfeafdd,
32'hbc06399a,
32'h3d40ac6e,
32'h3cd0e2bb,
32'hbc853210,
32'hbd983f76,
32'hbd496b40,
32'h3d502f0e,
32'h3d91af6b,
32'h3d7833ed,
32'h3cd2182a,
32'hbd552ad2,
32'hbc76a329,
32'h3c44d04d,
32'h3cc7b9df,
32'h3d45c0b1,
32'h3defac0f,
32'h3c97e13b,
32'hbdaeca1a,
32'hbdbe56ad,
32'hbb64e1e7,
32'hbbb97f32,
32'h3cfff37f,
32'hbd6d8a12,
32'h3d1d490f,
32'h3dc3f3b1,
32'h3d0139c6,
32'h3d8f4ff8,
32'hbde7273b,
32'h3b92ffc4,
32'h3d804f8e,
32'h3d76fd95,
32'hbd3efbf2,
32'hbdf28ae2,
32'hbd339291,
32'hbb4a12b9,
32'h3d4eae7d,
32'hbd50a4fa,
32'hbd13bf60,
32'hbdd830e5,
32'hbe0a80d5,
32'h3d37a054,
32'hbe807117,
32'h3c7dac56,
32'h3b7df32c,
32'hbd4b3eaf,
32'h3e690308,
32'hbc83a366,
32'hbd3ffd54,
32'h3d869650,
32'hbd90cf04,
32'hbd80d068,
32'hbe6318cb,
32'hbecb32a2,
32'hbdc2acc7,
32'h3efc807e,
32'hbd95adc5,
32'h3ecb6eaa,
32'hbdc9c41f,
32'hbe252c94,
32'h3e6fa464,
32'h3d9a8a50,
32'hbd9ee856,
32'hbe5ebef7,
32'h3d89ce9c,
32'h3c753fb1,
32'h3a377740,
32'hbcbb8528,
32'hbd8b8ce5,
32'hbcb314e3,
32'hbd2d64a3,
32'h3ccea804,
32'hbea4d45b,
32'h3a02f7ef,
32'hbdcc5c86,
32'hbd72c337,
32'h3e93c1c6,
32'hbc8c6c97,
32'h3d436e16,
32'h3bb6a15c,
32'h3e00566f,
32'hbdf9d67e,
32'hbe8ca517,
32'hbec52903,
32'hbe1e7abd,
32'h3eadff9c,
32'h3d5ba476,
32'h3ef860f7,
32'hbdad7db6,
32'hbca7fc55,
32'h3c896659,
32'h3d0ec077,
32'hbe78c042,
32'hbe272293,
32'h3dafab17,
32'hbd399399,
32'hbd5551ee,
32'h3e17dda8,
32'hbea6bdde,
32'h3d715739,
32'hbee97bf3,
32'h3dff22a2,
32'hbdf2253a,
32'hba438ce8,
32'hbd15004d,
32'hbcaf0eb4,
32'h3f15f7a7,
32'hbdee0490,
32'h3cb76c85,
32'hbd8bc901,
32'h3d8a6304,
32'hbdce70cb,
32'hbde2cbfc,
32'hbe7c8d92,
32'hbde426da,
32'hbc85b306,
32'hbe220d88,
32'h3f35a1bb,
32'hbdd03f8a,
32'hbd0324ff,
32'hbe4627be,
32'h3ce2ea3e,
32'hbdb0242f,
32'hbdc63419,
32'h3d0fe1ed,
32'hbd1e7c80,
32'hbc6fd95b,
32'h3f5a6ddb,
32'hbef100dd,
32'h3d6d8a07,
32'hbfaab745,
32'h3db3ea4b,
32'hbeba5f3c,
32'hbde19543,
32'hbc8f83dc,
32'h3ccb6438,
32'h3eced807,
32'hbfb29731,
32'hbd942f36,
32'h3f24991f,
32'h3dcfa2b6,
32'hbe6011dc,
32'h3d7ac763,
32'h3edb0c20,
32'hbd5406a4,
32'h3e5714bb,
32'hbe1d0c96,
32'h3fadfe02,
32'hbea49b83,
32'hbde9330a,
32'h3e635e57,
32'hbd6fbbc6,
32'hbf3b98a0,
32'h3db447a9,
32'hbd02797a,
32'hbd10e100,
32'h3f203210,
32'h3f665aca,
32'hbe2b1e3b,
32'h3cc06a2b,
32'hbf424982,
32'h3ecf796c,
32'hbf094c1c,
32'h3c6c0ad1,
32'hbd927697,
32'h3d39c5c4,
32'h3e53abe6,
32'hbf7d7d67,
32'h3efeb871,
32'h3f234ad3,
32'h3e05c132,
32'hbe621247,
32'h3d9b2162,
32'h3efd45aa,
32'hbd932696,
32'h3db56079,
32'hbd379224,
32'h3fb825fc,
32'h3e2f7f09,
32'hbd723f6d,
32'h3f1aa588,
32'h3c9bff53,
32'hbf235591,
32'hbde1ee53,
32'hbc7d4180,
32'hbd07b964,
32'h3ec5a59a,
32'h3e569601,
32'hbe8c911e,
32'hbea26887,
32'hbcd5bec8,
32'h3fbb0fd3,
32'hbdff3c61,
32'hbf04dbf9,
32'h3a5dc0ba,
32'h3d41f535,
32'h3fc1a3bd,
32'hbeda661c,
32'h3f24fb64,
32'hbf98efaf,
32'h3b0dcb95,
32'hbf3b4be2,
32'hbe3b7893,
32'hbf824c0d,
32'hbf500f89,
32'hbd9f5758,
32'h3f789205,
32'h3f2f238b,
32'h3e96b720,
32'hbcdbf473,
32'h3f8b1a95,
32'hbc263a56,
32'h3c722e09,
32'hbe9fb3b6,
32'hbcfe8b46,
32'h3a2af7ed,
32'h3e4447a3,
32'hbd2f63e9,
32'hbd192863,
32'hbe86df1d,
32'hbe6e31be,
32'h3f647b6e,
32'hbe3dd2eb,
32'hbea03808,
32'h3c693164,
32'hbd812780,
32'h3eca5a1f,
32'h3d526705,
32'h3f12bc8a,
32'hbf1225f4,
32'hbd002064,
32'hbe9fd82c,
32'hbd2430ce,
32'hbd9c0a98,
32'h3cfed3f9,
32'h3d8ff668,
32'h3f5065e6,
32'h3ef67f44,
32'hbe17c9c4,
32'hbd4613af,
32'h3e0134af,
32'hbd39fb5c,
32'hbe3fad7c,
32'h3e85b4b4,
32'h3d169425,
32'hbce0adc7,
32'hbe62ddc9,
32'h3e087cee,
32'hbd8e4f7a,
32'hbf063dd1,
32'h3f204b5d,
32'h3fdc0a23,
32'hbe1eb693,
32'h3ea618a1,
32'h3d06b77f,
32'hbcd0e3f2,
32'h3f2c5add,
32'hbe142d0a,
32'h3e6c5d3d,
32'hbeb74f51,
32'h3fa1acef,
32'hbf7d1c54,
32'hbf23313e,
32'h3e488dde,
32'hbeda2984,
32'hbe808795,
32'h3e80d598,
32'h3ef2d9ae,
32'h3cb58443,
32'hbd140ef8,
32'h3f0a052d,
32'hbda3a31c,
32'h3f5bdaca,
32'hbda07e17,
32'hbe3b4373,
32'hbdf9097c,
32'hbe948b43,
32'h3e49cef8,
32'hbd5989a0,
32'hbe068329,
32'hbe7b3a13,
32'hbe90f5fa,
32'hbcf97785,
32'h3e82318e,
32'hbcaedbc0,
32'h3dc71e63,
32'h3e7f124e,
32'hbeeebb93,
32'hbe268e87,
32'hbdf4df20,
32'h3f929f65,
32'hbdffb5bc,
32'hbe75317a,
32'hbe63b306,
32'hbcc1eb7a,
32'hbe3bd6a0,
32'hbef8eee8,
32'h3f2c28c8,
32'hbddb38e1,
32'h3cc444ad,
32'hbe6dfed9,
32'hbd7e5178,
32'hbd5f1b8f,
32'h3f175e08,
32'hbec1ee4b,
32'hbe8a3000,
32'h3e029df0,
32'h3d3d9e0d,
32'hbe5bb66c,
32'h3cc79bcf,
32'hbec8c766,
32'hbf0b5b43,
32'h3eb801de,
32'hbe22feb6,
32'h3c90c3d5,
32'hbcb501a1,
32'h3f3d56e0,
32'hbe649e49,
32'h3e7dfbe9,
32'hbf031d97,
32'h3fbdf509,
32'hbf81ad7f,
32'hbfc836c4,
32'hbfa49672,
32'hbeb29eee,
32'h3e264118,
32'hbe8600af,
32'h3f92ee8b,
32'h3d521d68,
32'hbea9f242,
32'h3c872d6b,
32'h3d76e0c0,
32'h3e1b89e6,
32'h3f0a03fe,
32'hbfc5a451,
32'hbdd576fa,
32'h3fa301ba,
32'h3e4be5fd,
32'h3dfdde95,
32'h3d3c7b85,
32'hbf07945a,
32'hbe41aefe,
32'h3f8d6131,
32'hbf78fdd3,
32'hbc6b4ba8,
32'h3c4cb29a,
32'h3ef3fe41,
32'h3f146511,
32'h3fb5837d,
32'hbf91ef7e,
32'h3f7ee21d,
32'hbd91adef,
32'hbf5d750d,
32'hbf9913cf,
32'hbeb44575,
32'h3e9fab9f,
32'hbf9b5f44,
32'h3ec728ee,
32'h3f2681d1,
32'h3d82fda5,
32'h3e283f85,
32'h3d4a8081,
32'h3f86423e,
32'hbe5af2f8,
32'hbe972fb9,
32'hbcf44296,
32'h3f642f92,
32'h3e52e8c3,
32'h3e80530d,
32'h3e2282e0,
32'hbe1e8525,
32'h3e893165,
32'h3de96f30,
32'hbe111253,
32'hbdc24e07,
32'hbda1df5a,
32'h3f7a37e6,
32'hbc5873d2,
32'h3ebf1e2a,
32'hbf544356,
32'h3f629f28,
32'hbdc8b186,
32'hbd989ac7,
32'hbf8a5b77,
32'hbe5b08ce,
32'h3e002a89,
32'h3ea665ea,
32'h3ecfa7e8,
32'hbe26c362,
32'hbbf2ee9d,
32'h3e0fc58d,
32'h3b8acd42,
32'hbe67d6e7,
32'h3e03807a,
32'h3d831c95,
32'h3c04acd0,
32'h3e379753,
32'hbea3f7ff,
32'hbd8d32ae,
32'h3d2326e3,
32'hbd90fcbe,
32'h3e8e7ae9,
32'hbe550c12,
32'hbf36b2ce,
32'hbd091962,
32'hb9878c51,
32'h3f902441,
32'hbe14d20c,
32'hbe322205,
32'hbfdabe2c,
32'h3ef9bfb4,
32'h3dcc9dfb,
32'h3ddf8d2d,
32'hbf0e2c72,
32'hbe7e159a,
32'hbeaffd91,
32'h3f94c702,
32'h3f09e808,
32'hbdc1932b,
32'hbd7d0f9a,
32'hbeefc6c7,
32'h3f52c0b1,
32'hbe63f5ae,
32'hbcee0475,
32'h3d5c0e69,
32'hbc54418d,
32'h3cbb47fc,
32'h3d9c438d,
32'h3d2bcc3e,
32'h3e869704,
32'hbeef4e2a,
32'hbe42202a,
32'h3f1e48f1,
32'h3d026092,
32'h3dcf621c,
32'hbd223d72,
32'h3f5696a9,
32'h3d42c83b,
32'h3d9cf061,
32'hbdde3c17,
32'hbd4572ce,
32'h3cef5f70,
32'hbf0f5a12,
32'h3ee9d315,
32'hbdce1dac,
32'hbe0c2246,
32'hbe91974c,
32'h3a8a9fd5,
32'h3d0acc95,
32'h3d7b766e,
32'hbdbc2e36,
32'h3d2d8e49,
32'hbda75c35,
32'h3de67526,
32'hbc9e1e14,
32'hbc3ac621,
32'h3c235d1c,
32'h3c685a7e,
32'hbc8857c0,
32'h3ea06c7d,
32'hbd9a396e,
32'hbdf21e70,
32'h3f0b03b6,
32'hbd130b3f,
32'h3e11b382,
32'hbd441b70,
32'h3f534eef,
32'h3c4c380c,
32'hbd99004a,
32'hbe8e95ad,
32'hbce296d3,
32'hbde7d826,
32'hbeca74fb,
32'hbed3dc13,
32'hbe4ed6f1,
32'h3d3c3702,
32'h3ecd9b2e,
32'h3e87faeb,
32'h3a90d295,
32'hbd2cd00f,
32'h3d51d9a1,
32'hbd6e4749,
32'hbd62398a,
32'hbb188f7f,
32'h3da43022,
32'h3db11107,
32'hbc22c542,
32'hbc14e9de,
32'hbce738f9,
32'h3ee50435,
32'hbeca336b,
32'hbe4b48b2,
32'hbd97d138,
32'h3c0f2e85,
32'h3cef3ce8,
32'hbc13c2f7,
32'h3f276d55,
32'hbe283f7b,
32'hbe40544b,
32'hbc8c8ac9,
32'h3d6f987d,
32'hbd9eb86c,
32'hbe41d094,
32'h3e138c36,
32'hbd5b0f6b,
32'h3e0575b4,
32'h3e40d756,
32'h3d1ba13f,
32'h3deccc60,
32'hba2748a5,
32'hbe401661,
32'h3cb38dc0,
32'hbc5ab015,
32'hbce1e069,
32'h3d84cfde,
32'h3d194051,
32'h3dc670f5,
32'hbbb4e4f5,
32'hbe0ab35e,
32'h3ec9f361,
32'hbe8b46c4,
32'hbec78f00,
32'hbe79b9f8,
32'h3e015956,
32'h3d99eef6,
32'hbddb0d26,
32'h3f617290,
32'h3d0aba36,
32'hbe426c60,
32'h3d41a358,
32'h3d88b836,
32'hbd06b80b,
32'hbe8f9ce7,
32'h3e729ce1,
32'hbdbf72f1,
32'h3d04cac3,
32'h3ded1eb7,
32'h3e2e74bc,
32'h3e8ad846,
32'hbd0d1597,
32'hbe4697ed,
32'hbda2aed2,
32'hbd47bebf,
32'hbe3ba611,
32'hbd5fc76d,
32'h3d6fb2c4,
32'hbb90fc5f,
32'h3d9b87cb,
32'h3cc8f19e,
32'hbd938372,
32'hbd15dd60,
32'h3ce0ded6,
32'hbd862fa2,
32'hbc89d264,
32'hbde36f48,
32'h3d106e7d,
32'h3e07d0f0,
32'hbd4e663b,
32'h3d184338,
32'hbd9b01dc,
32'h3cc1e375,
32'hbdedd5fa,
32'hbdc86f74,
32'hbd0f3ea9,
32'hbe17b54a,
32'h3dd163e5,
32'hbcdf5700,
32'h3d0f00bd,
32'h3c802cc5,
32'h3c908496,
32'h3d3d8eee,
32'hbbc486b7,
32'hbcc7f6b3,
32'hbd3439bf,
32'hbd464d6e,
32'h3ba202d5,
32'h3dc11771,
32'h3d81e00a,
32'hbc47072a,
32'h3c95d909,
32'h3c609c07,
32'h3d1d14f6,
32'hbc9d51a2,
32'h3d805157,
32'h3dc46d09,
32'hbd3c8719,
32'hbd7c49db,
32'hbc2cab23,
32'hbdb66cf7,
32'hbd44f892,
32'hbcc4b4e3,
32'h3d263d3b,
32'h3c1c39a7,
32'h3c94baad,
32'h3c9fc499,
32'hbcc0a731,
32'h3d6c1ae6,
32'hbd8b2d32,
32'hbb053c82,
32'h3c7bf5d3,
32'h3d7abd38,
32'hbdb8a69a,
32'hbc959660,
32'hbd8868be,
32'h3cb3c4a0,
32'h3cdc4f19,
32'h3d78b110,
32'h3cd6c1e9,
32'hbd2f4b5d,
32'hbd06e9b9,
32'hbc74ee71,
32'hbd8a5e81,
32'h3cfff487,
32'h3d56f591,
32'h3dd95ac1,
32'h3cd72606,
32'h3d249554,
32'h3c57d851,
32'hbd02f9be,
32'h3d16f4e1,
32'hbde9aff5,
32'h3d9733fb,
32'h3d967e70,
32'hbd5a2a51,
32'h3c90bebd,
32'hbcb50bf0,
32'hbba89d40,
32'hbcc2eb09,
32'hbdbc693b,
32'hbc1e9c44,
32'h3cbb4405,
32'h3da2c262,
32'hbd17b4bb,
32'hbd3422e5,
32'h3d151894,
32'h3d89f7de,
32'h3dc68861,
32'h3c74221f,
32'h3c5df82c,
32'h3d2de35b,
32'hbc5139b2,
32'h3d15342c,
32'hbdb8f14c,
32'hbd73a105,
32'hbd83238f,
32'hbcb5c580,
32'hbd97a97c,
32'hbce9d2dc,
32'hbd8854cc,
32'hbcef9450,
32'hbc41f6bd,
32'hbd048e47,
32'hbdc6561c,
32'h3da2fafe,
32'hbbe4592b,
32'h3bb6ddf8,
32'h3db17857,
32'hbd4f7dc1,
32'h3db076ff,
32'h3ca280ba,
32'h3ae90beb,
32'hbd061f37,
32'h3da346bc,
32'h3d08c136,
32'hbb59cf1e,
32'hbd07647f,
32'h3d2cf0f0,
32'hba3c8e3d,
32'h3cc74005,
32'h3d24a083,
32'hba1cb26c,
32'h3d3960c8,
32'hbd14b225,
32'hbd47584e,
32'h3da72ef6,
32'hbc3d6ac9,
32'hbce79520,
32'hbce4307b,
32'h3d7f13bd,
32'h3cee6fdb,
32'hbbe34285,
32'hbd0e7999,
32'hbb96ad3d,
32'h3d9c1275,
32'hbbd4fd7c,
32'hbca12e59,
32'h3d5228ac,
32'hbce862ae,
32'hbca54c89,
32'hbb9c27af,
32'hbcd563ca,
32'h3da87712,
32'hbd739588,
32'hbba03387,
32'h3c866843,
32'h3dbc22cd,
32'hbd258a29,
32'hbd43f940,
32'hbd809ea2,
32'h3d70c2c1,
32'h3ac7aac6,
32'hbd181ffe,
32'h3d2d1327,
32'h3d9a7c78,
32'hbc8204cf,
32'hbd5dccf4,
32'h3d7a3043,
32'hbcdbc1c7,
32'hbc5b7959,
32'hbd191039,
32'hbd5cf464,
32'h3c4e7a60,
32'h3b3dbc14,
32'hbc10d58b,
32'hbdb8b862,
32'hbde5f8e4,
32'h3cf76c6e,
32'h3d217abc,
32'hbde44274,
32'h3d1b8561,
32'h3d233524,
32'h3d90f9f4,
32'hbc613db9,
32'hbd85729e,
32'hbc7ccc03,
32'hbd192367,
32'h3d047dfd,
32'h3c4948c8,
32'h3d7c6175,
32'hbd084ce0,
32'h3c4c787a,
32'h3c8e4aa0,
32'h3d6a131c,
32'h3dacc44f,
32'hbc6daec2,
32'hbd220def,
32'hbcf08f0e,
32'h3cffd35b,
32'h3d30aa84,
32'h3d3dba51,
32'h3bd07790,
32'hbd1fe665,
32'hbdb35900,
32'hbd8f0c0a,
32'h3db75ae8,
32'hbd3064c0,
32'hbdafd22d,
32'hbd512f33,
32'hb9922f2d,
32'h3b316483,
32'hbd7b5a0d,
32'h3cdc0963,
32'hbd79b5ab,
32'hbceaed86,
32'hbd8d87d5,
32'hbcbf434c,
32'h3c8f57d1,
32'h3d0af598,
32'hbbe03b52,
32'hbccd33d0,
32'h3c9e6312,
32'h3d17cbe3,
32'hbcfe6308,
32'h3d98b785,
32'h3dba9511,
32'h3c4411fb,
32'h3ce666f2,
32'h3ce4aba2,
32'h3d964d88,
32'h3af9ffe2,
32'h3ce3bf8f,
32'hbb854cac,
32'hbd905661,
32'h3d91f96f,
32'hbddeb4ab,
32'h3d5b455e,
32'hbd71732f,
32'hbd808650,
32'h3b60d238,
32'hbcf5583e,
32'h3c1bc65d,
32'h3d0dcd16,
32'h3d43c752,
32'h3cda0264,
32'hbdc6c5fa,
32'h3c16983e,
32'h3b4d1ff0,
32'h3ea2aee0,
32'h3d173404,
32'hbdb3eefc,
32'h3d19c02f,
32'h3e76e75d,
32'hbc1f3e6c,
32'hbcbd843c,
32'h3c8f19e8,
32'h3cf01b75,
32'h3ecf3f24,
32'h3d104292,
32'h3cc4cb75,
32'hbea051a6,
32'hbccf47fc,
32'hbd895ca1,
32'hbdf9f974,
32'hbeac2cfb,
32'h3d86025c,
32'h3cdf3f71,
32'h3ccadb0d,
32'h3dba3e06,
32'h3a2c7842,
32'h3d8ebbdf,
32'h3d2bf604,
32'h3bd2fd65,
32'hbd221c33,
32'hbecbeacc,
32'h3c7883b9,
32'hbc937cfa,
32'hbbd57d8b,
32'h3e890736,
32'hbd211aa2,
32'h3dd93c10,
32'h3b95a6e5,
32'h3e522635,
32'hbce59c77,
32'hbd324158,
32'hbcefae16,
32'h3cf8fa5a,
32'h3ebae96a,
32'hbc376965,
32'hbc7b7b3a,
32'hbeb7f063,
32'hbd42bc73,
32'h3c9335eb,
32'hbded251d,
32'hbe7405da,
32'hbc9e7eee,
32'h3de2946c,
32'hbc6a6b19,
32'h3bbc4e8a,
32'h3dab5e08,
32'hbd907973,
32'h3d75c6c0,
32'h3b4f06d0,
32'hbcabb71c,
32'hbebaf6cf,
32'hbce101e4,
32'hbd16e874,
32'h3da4c9a1,
32'hbd8b30ab,
32'hbd9775c2,
32'h3d2aa77b,
32'hbd0de78b,
32'hbdff5b70,
32'hbdda7093,
32'h3bd085da,
32'hbd5b6388,
32'hbd06c58e,
32'h3e2cd14c,
32'h3e4b42c7,
32'h3ddc9d54,
32'hbd420067,
32'h3df1d29c,
32'hbd28fda7,
32'hbd758fce,
32'hbe3b4ba4,
32'h3cc9f6b1,
32'h3dc8b567,
32'h3d3668f3,
32'hbd4a83bd,
32'h3e06e983,
32'hbdc80ec9,
32'h3e2ce6f2,
32'hbd32243c,
32'hbcb30c73,
32'hbe5ce313,
32'h3dbf9b16,
32'h3ddb4fb7,
32'h3eb37a9e,
32'hbdf7c278,
32'hbdc64b0b,
32'h3db3b267,
32'hbd9e5829,
32'hbde1e8be,
32'hbd9c3fc6,
32'hbdc753e4,
32'hbd439800,
32'hbdc959e3,
32'h3e9e0351,
32'h3eb76923,
32'h3e0e65c8,
32'hbe3bf327,
32'h3e84748a,
32'hbe30d792,
32'hbe601bb0,
32'hbe55c0a5,
32'hbd2450ac,
32'h3ea72040,
32'hbdc1ac96,
32'h3f12b50e,
32'h3d460dba,
32'hbd5a8674,
32'h3e1a7d72,
32'hbc898efc,
32'hbe3744a1,
32'hbec970b8,
32'h3d94a4ad,
32'h3e03d517,
32'h3e6e5eb0,
32'hbe94a8bd,
32'hbe2bf1f9,
32'h3d308a92,
32'h3ef04a4b,
32'h3f3c1e23,
32'hbe6503f3,
32'hbcccb03a,
32'h3d2ec69e,
32'hbd0d0b57,
32'h3e3a6afc,
32'h3f732f3a,
32'h3ea0fa29,
32'hbcd30838,
32'h3ed17424,
32'hbdc29f8b,
32'hbe948cdb,
32'hbebfc8e9,
32'hbde65c39,
32'h3e98d7eb,
32'hbe799798,
32'h3f28ca07,
32'h3e01203d,
32'hbc87d80c,
32'hba524842,
32'hbd3c2eac,
32'h3e1eb135,
32'hbe950dce,
32'hbce06798,
32'h3cfd7477,
32'h3e7c29cb,
32'h3e7fb8f1,
32'hbf0b9a50,
32'hbf45ea22,
32'h3f291fc2,
32'h3eb22455,
32'h3e2e2404,
32'h3f50cf81,
32'hbab66d84,
32'h3dd89532,
32'h3f53aba7,
32'h3e09c341,
32'h3db23521,
32'hbbd683bf,
32'h3fe7ab0b,
32'hbe968c01,
32'hbe2c84d6,
32'h3d57d41b,
32'hbe2602af,
32'hbeefd3ee,
32'hbe88f1d7,
32'h3f42f8de,
32'h3f243984,
32'hbdc60c0d,
32'hbe125d1c,
32'hbe69af67,
32'h3e9ca806,
32'hbe37f019,
32'hbb19a91f,
32'hbe09cf29,
32'hbd665f6a,
32'hbff25931,
32'h3ec4c646,
32'hbf15a0e2,
32'h3f3851e7,
32'hbe350975,
32'h3ef240a8,
32'h3e949e9e,
32'hbd114798,
32'h3d6fa2cb,
32'h3f9f2dd3,
32'h3ece4e88,
32'h3edf2f0a,
32'hbf01b839,
32'h3fd22286,
32'hbe87fae6,
32'hbe805b6e,
32'h3ec33d95,
32'hbe18b57b,
32'hbf0cf407,
32'hbf27f07e,
32'h3fee8f9d,
32'h3e4512ef,
32'hbb804f0f,
32'hbf100cae,
32'hbeba8f72,
32'h3f6b8261,
32'h3e6e7f6d,
32'h3db75468,
32'hbe235dc2,
32'h3e649fb5,
32'hbe402c89,
32'hbf0de109,
32'hbf7cde25,
32'h3e3dc1fc,
32'h3f83f7e4,
32'h3d3d9c3a,
32'h3f0cea74,
32'hbdcc674f,
32'h3c7a40e9,
32'h3f99487d,
32'hbbf8edae,
32'h3f3f86eb,
32'hbf2276dd,
32'h3f374198,
32'hbf06b05b,
32'hbf3009c3,
32'h3e78bc64,
32'hbf5cd049,
32'h3db782ff,
32'hbea22263,
32'h3fd30e98,
32'h3f12a27c,
32'hbd168aee,
32'hbe6a5564,
32'hbe924031,
32'h3f8154ff,
32'h3ed7652e,
32'hbc9122c6,
32'hbeb311dd,
32'h3f29b8d1,
32'hbf62e24c,
32'hbe3f3fef,
32'hbf0f0079,
32'h3f5efdc3,
32'h3f6b66e2,
32'hbd90eb10,
32'h3f64a6d8,
32'hbd758d92,
32'hbd879329,
32'h3f6fa6de,
32'hbd940b7a,
32'hbd327234,
32'hbf54d851,
32'h3dbce68b,
32'hbfbe53b3,
32'hbfcc76a4,
32'h3e1e1845,
32'hbf69e105,
32'hbd4f8ad8,
32'h3e03f763,
32'h3fd0bc12,
32'h3eca80ab,
32'hbe00ca95,
32'h3e85c731,
32'hbf139db0,
32'h3f916c50,
32'h3f3e67dd,
32'hbed0797a,
32'hbe2de032,
32'h3fc42ab8,
32'h3cc56b15,
32'hbd5b72d3,
32'hbfcfbad6,
32'h3e875bc6,
32'h3d67e7b5,
32'hbdff4635,
32'h3e2a5f36,
32'hbdb2654d,
32'hbd3abf0d,
32'h3fe64c3f,
32'hbe5a27fa,
32'h3d34df96,
32'h3eca607c,
32'h3eacc030,
32'hbf8a13ab,
32'hbfd86f9f,
32'hbf0905d9,
32'hbf10b10b,
32'h3ec6d6b3,
32'hbfc3d526,
32'h402a8ee6,
32'hbece661a,
32'hbd946f7d,
32'h3f77993c,
32'hbe58743d,
32'hbdd08954,
32'h3efece87,
32'hbec56fa1,
32'hbeb9ed17,
32'h3ea3121f,
32'hbee615e9,
32'hbe84a576,
32'h3e1cf80f,
32'h3e6ba461,
32'hbc831132,
32'h3db245b5,
32'h3f627538,
32'h3d9b2e56,
32'hbdcb5e3f,
32'h3f7b3f15,
32'h3ea5d768,
32'h3ea10b76,
32'hbe83ec7a,
32'h3f95b71b,
32'hbf82cd27,
32'hbfd5e681,
32'hbf05cb49,
32'hbf1faa0a,
32'h3b25dd64,
32'hbfb04bb7,
32'h40025f61,
32'h3f01ad4b,
32'hbcfc529a,
32'h3d5216ed,
32'h3b1da826,
32'h3f80c824,
32'h3f07ec2b,
32'hbef71a17,
32'hbf4b8d79,
32'hbf266e2a,
32'hbfb4cb8b,
32'hbeadef7e,
32'h3d9a6c45,
32'hbf1a03cc,
32'h3e269b5d,
32'hbf3831b5,
32'h3eb482f1,
32'hbd8893e0,
32'hbd05e164,
32'h3f07fbb5,
32'hbeb8fce4,
32'h3f3920a0,
32'h3e066ae1,
32'h3e415c56,
32'hbfa1149c,
32'hbfd8864a,
32'h3f5fa696,
32'hbf9897bc,
32'hbe528484,
32'hbde617ff,
32'h3f915fe5,
32'h3f18de29,
32'hbf021a00,
32'hbe69cda4,
32'hbeb9d308,
32'h3f0d34a0,
32'h3f2bafe1,
32'hbfc44d45,
32'hbf0c7f76,
32'hbf808331,
32'hbfb5f3c8,
32'hbe0afe9e,
32'h3ed3c293,
32'hbf719877,
32'h3e97c5f2,
32'hbf17b2a8,
32'h3ea5ecee,
32'hbd2ae533,
32'hbd89a91f,
32'hbf216301,
32'hbf7a059e,
32'h3f58bc4e,
32'h3f74576e,
32'h3ebd28e1,
32'hbf2f5921,
32'hbf8431db,
32'hbd6d06ff,
32'hbeafc825,
32'hbe1cb029,
32'h3dbb1e1d,
32'h3f180ff1,
32'h3ee478fb,
32'hbf5939cf,
32'h3df335ae,
32'h3dd85327,
32'h3f2a6572,
32'h3e736341,
32'hbffa1572,
32'hbf2cc308,
32'hbfa0cc0c,
32'hbfc244f2,
32'hbe47bf3a,
32'h3e67651c,
32'hbf73085f,
32'h3e9254e7,
32'h3e87457a,
32'h3f76e245,
32'hbd891489,
32'hbc113fea,
32'hbd4179c9,
32'hbf2d83b9,
32'h3e918926,
32'h3ec43201,
32'hbd9c4252,
32'hbd23f815,
32'hbfceaacd,
32'h3ceed741,
32'hbe909848,
32'h3e306d99,
32'h3ea3e61a,
32'h3e426dd8,
32'hbeb2cfc4,
32'hbf14c5fe,
32'hbebb8fe8,
32'h3d804995,
32'h3f6715df,
32'h3e33ad61,
32'hbfd36023,
32'hbf2f2903,
32'hbfb9be1e,
32'hbf72c9e3,
32'hbf1ba3ef,
32'hbedf246a,
32'hbf78ce87,
32'hbeb86bce,
32'hbe6c5292,
32'hbf904489,
32'hbe0be2a2,
32'h3d3d5d5a,
32'hbb22effa,
32'hbef54c09,
32'h3d7e6fd8,
32'hbeb59d93,
32'hbed76afe,
32'hbeb44ff0,
32'hbf8ce435,
32'h3e1ec56f,
32'hbf86119c,
32'h3ec75d74,
32'h3edc368c,
32'h3f7d47a6,
32'hbeb28a3b,
32'hbefc9b2e,
32'hbf3197fc,
32'h3f296662,
32'h3f062e54,
32'hbe2d55a4,
32'hbfc05ea9,
32'hbebd578b,
32'hbf96028d,
32'hbfd1ddab,
32'hbf283de7,
32'h3ef76fd1,
32'hbff15fd3,
32'h3e33382f,
32'h3cb10b2a,
32'hbfe5785a,
32'h3d2421e3,
32'hbd4e714f,
32'hbe5b1e4c,
32'hbf54159a,
32'hbe01311c,
32'hbf0a5ad7,
32'hbfd2693b,
32'hbf3783ec,
32'hbfa43623,
32'hbf3cacfd,
32'hbf7d3253,
32'h3f174b1b,
32'h3e743da2,
32'h3f5b4773,
32'hbeaae2fe,
32'hbdacc42b,
32'hbe90a486,
32'h3f9b0036,
32'h3e6dfc68,
32'hbf18137b,
32'h3d091fbf,
32'hbdc1fe76,
32'hbeaa197f,
32'hbff75b0d,
32'hbee1bf95,
32'h3ecb2b5a,
32'hbf98ffbc,
32'hbf27bbed,
32'hbe19e9dc,
32'hbf5f6043,
32'h3d22e4ce,
32'hbd412c48,
32'h3efee763,
32'hbf9b2836,
32'hbd75b6c1,
32'hbf655461,
32'hbfd30f7b,
32'hbed30f9b,
32'hbf9ff794,
32'hbe6810c2,
32'hbf924ca5,
32'h3f0a6906,
32'h3f73544d,
32'h3f90488e,
32'hbee19ecf,
32'h3d3700bd,
32'hbf081774,
32'h3f453746,
32'hbe92ccc2,
32'hbf29ed3b,
32'h3e91ff9a,
32'hbd39da38,
32'hbf312c01,
32'hbee27dc4,
32'hbeb3ca87,
32'h3e874465,
32'hbf00bcef,
32'hbeae1ff9,
32'h3f2e1a94,
32'h3de65fb7,
32'h3c36ded2,
32'hbdf41ee7,
32'hbe490b9f,
32'hbf31428b,
32'hbdc323a7,
32'hbe7ead0f,
32'hbfe53b81,
32'hbbc44789,
32'hbfa59979,
32'h3dde7e1c,
32'h3f0f06de,
32'h3f13831e,
32'hbd82d8ee,
32'h3f21fd4c,
32'h3ed31c71,
32'h3d002ba1,
32'hbd8a619f,
32'h3ef60d47,
32'hbe868d6e,
32'hbe7ccdde,
32'h3e36731d,
32'hbcf46e5d,
32'hbe58d89f,
32'h3e5e3ff4,
32'hbe8ff87f,
32'hbe2467b5,
32'h3e85875c,
32'h3d20cf30,
32'h3f17fe2a,
32'h3e03fa5a,
32'hbd63bc63,
32'h3dc75926,
32'h3dad88f1,
32'h3f8dd088,
32'h3f0f8b3a,
32'hbf6e7133,
32'h3f5e6351,
32'h3ec5f982,
32'hbf1f38fe,
32'h3e2245ed,
32'h3f37ae89,
32'hbe32dc6e,
32'h3e5e3321,
32'h3ea16d77,
32'h3f0f651b,
32'h3c76eb31,
32'hbca5d81e,
32'h3ec8c3c6,
32'h3e5a03bd,
32'hbe3d0398,
32'h3db6415e,
32'hbba4e492,
32'hbda64efb,
32'h3e3a0188,
32'hbe7bfef9,
32'h3eab90e6,
32'h3e6de6dc,
32'h3e92a26b,
32'hbdc3704f,
32'h3eebf841,
32'h3d113498,
32'hbc26367b,
32'h3e1bda2a,
32'h3d398221,
32'h3d1cc698,
32'hbf273df5,
32'hbd74081a,
32'h3f2e75ab,
32'hbdb2c389,
32'h3eaa2672,
32'h3e46385e,
32'hbd804f37,
32'h3dd9b1c7,
32'h3f1b28fe,
32'h3e053cfb,
32'h3c9946f2,
32'hbecfa68c,
32'h3ea19092,
32'hbdb3c310,
32'h3e96583a,
32'h3c6e132e,
32'h3b4d17ef,
32'h3f7e2986,
32'h3d86895b,
32'hbdd41da0,
32'hbf12547d,
32'h3f49d84a,
32'h3eef1582,
32'h3f5211e3,
32'hbc5b696e,
32'hbca5baf0,
32'h3d3066c4,
32'h3e0a7c76,
32'h3eb85740,
32'h3f797020,
32'hbf922776,
32'h3e7eb644,
32'hbd9c8421,
32'hbe6300da,
32'hbed18b79,
32'hbe3aa58b,
32'h3dc161b6,
32'hbd4a3525,
32'h3e175515,
32'h3edc0d69,
32'h3d4576b5,
32'hbe7ccb84,
32'hbd9c8590,
32'h3f84b3b6,
32'hbe3cc699,
32'h3c120a17,
32'hbd7bb245,
32'hba3bb392,
32'hbdaa09e5,
32'hbbe36f89,
32'hbe503d15,
32'h3f572613,
32'hbb9c8235,
32'h3f44e0ce,
32'hbd143e6b,
32'h3c8833de,
32'hbd1002bc,
32'h3dcf314f,
32'h3ecc40ce,
32'h3c933036,
32'hbe8508bc,
32'hbd7523db,
32'h3d4c68f7,
32'hbd5f85bb,
32'hbc785e10,
32'hbca2e83c,
32'hbe9fbf7e,
32'hbd98e760,
32'hbe9f3ffe,
32'h3e833e91,
32'h3bf31a1f,
32'h3f106931,
32'hbd25ebd1,
32'h3f1a28da,
32'hbc8888c9,
32'h3daa758c,
32'hbcc05dcb,
32'hbcec7826,
32'h3b703f0a,
32'hba829f57,
32'hbe8daa3b,
32'h3f5ec4bf,
32'h3d29dac8,
32'h3f444363,
32'h3c8b9f65,
32'hbdc2698f,
32'hbdb0da3e,
32'hbe99591d,
32'h3f435775,
32'h3df38f43,
32'h3d8537ae,
32'h3dddbf80,
32'h3c3180a5,
32'hbdbcac75,
32'hbc967dbe,
32'hbad7a608,
32'hbe2feb17,
32'hbe5a416c,
32'hbf5e4a4a,
32'h3e3d1176,
32'hbda282ed,
32'h3f4625f7,
32'hbda1d70f,
32'h3f1f9ab0,
32'hbe893379,
32'hbdb4fbaf,
32'h3cdc8a6a,
32'h3d844527,
32'h3d98e838,
32'hbdb8089c,
32'hbce3418a,
32'h3d7607b4,
32'h3ddd8afc,
32'hbc9a08e9,
32'hbde0aaf7,
32'h3dba9b64,
32'hbca892d4,
32'hbc086482,
32'h3cd51a0a,
32'hbcdc8510,
32'h3d215cb3,
32'h3d8c9cde,
32'h3d4cf247,
32'h3be3dd5f,
32'hbdc13550,
32'hbd00fd83,
32'hbd5c4f57,
32'h3c12f167,
32'h3cca4da5,
32'hbcbfa792,
32'h3b13df14,
32'hbbe0885e,
32'h3dd5d65e,
32'h3cac83b3,
32'hbbb928fc,
32'h3cce5b7e,
32'h3d105c0f,
32'hbbbc6dbc,
32'h3d4f8d5c,
32'hbbc1e88e,
32'hbd2aa0a4,
32'h3c6dfe54,
32'hbcf7e19a,
32'hbd47ee8f,
32'hbd3d2383,
32'hbd3ce022,
32'h3d7c3a69,
32'h3dacc200,
32'h3c476567,
32'h3cf1ca11,
32'hbd3c2278,
32'h3daf2c3b,
32'hbda9afeb,
32'h3c73f74f,
32'h3b9e26b3,
32'h3db73dd1,
32'h3d524a0d,
32'h3c16ed36,
32'h3d64364f,
32'h3dcd66eb,
32'h3dabd93a,
32'hbc406728,
32'h3d84a8ab,
32'hbdcf0f75,
32'h3d690e81,
32'hbdcb6f6f,
32'h3d44df7e,
32'h3d415e50,
32'hbd4e6de1,
32'h3ce5ec2d,
32'h3969181c,
32'hbc07c03a,
32'h3cd60cf5,
32'h3db380e2,
32'hbc6e7fff,
32'h3d187320,
32'h3c7d03bb,
32'h3d06f677,
32'h3d0fecf3,
32'hbdd48bca,
32'hbd80b170,
32'h3da9feff,
32'h3d4f6a9b,
32'hbcd9f062,
32'hbc21bc16,
32'h3d348e68,
32'h3cc739c4,
32'h3b4182f0,
32'h3c203c09,
32'h3c8e58c8,
32'hbd0abd24,
32'h3befc81d,
32'h3d8d5c85,
32'h3d32499b,
32'h3d22ac14,
32'h3c56394f,
32'h3d805a31,
32'h3d4ae6ec,
32'h3dda8007,
32'h3d87b8d6,
32'hbc9cbb74,
32'h3caa253d,
32'hbd1e0e86,
32'hbd0c2fb7,
32'h3d8bc46a,
32'h3d28fe97,
32'h3d988be4,
32'h3d45e586,
32'h3d612e66,
32'hbc9f861d,
32'h3cf624cb,
32'h3d9094cc,
32'hbd8b41ef,
32'h3a814994,
32'hbccd8c07,
32'h3d1d8c56,
32'h3c1529d5,
32'h3d5fa168,
32'h3d61a280,
32'hbd7f3483,
32'hbc13c3a9,
32'h3d8d62e9,
32'hbcb15b8b,
32'hbd94a5c6,
32'h3d331129,
32'h3ee8bced,
32'h3a9fa98b,
32'h3db98efa,
32'h3c598394,
32'h3b8cafe2,
32'h3d955ff8,
32'hbd1ba75a,
32'hbe2b2145,
32'h3d65ca6f,
32'h3f5467a6,
32'h3d8fd9ad,
32'hbc39b8d0,
32'h3d1208ab,
32'h3e056bdf,
32'h3d8f77c2,
32'h3f214827,
32'h3d88a1bc,
32'hbcb7d378,
32'h3dbd2a3c,
32'h3bb6d1c1,
32'hbe2f0cea,
32'hbef73fce,
32'hbf328225,
32'hbf5603d5,
32'hbe3ca2be,
32'h3c9b28c5,
32'h3e113e77,
32'hbd134e8e,
32'h3d0cdd4f,
32'hbe9e9ce0,
32'h3f074059,
32'hbdc62ff4,
32'h3cb6aaa7,
32'h3dd6b7e6,
32'h3d9c4712,
32'h3cff5509,
32'hbdede00e,
32'h3f136ecc,
32'h3da7647e,
32'h3f33c5aa,
32'hbd6ce923,
32'hbcf3f725,
32'h3ea1220b,
32'h3e8edd8d,
32'hbd17fee0,
32'hbd6306ac,
32'hbd882c25,
32'hbecc616f,
32'hbe5508dd,
32'hbf2c15f8,
32'hbe52dca0,
32'h3d117996,
32'hbf419788,
32'hbebb29cd,
32'hbc2e9454,
32'h3d25e6a3,
32'h3f243deb,
32'h3cb7688f,
32'h3d575768,
32'hbf76a587,
32'hbd6b1b15,
32'hbe206339,
32'h3e4e561e,
32'h3ec60633,
32'h3d5e1790,
32'h3e098d4e,
32'hbd85168e,
32'h3e85a0d7,
32'h3af67787,
32'hbd9e306d,
32'h3d5e93ed,
32'hbd92e128,
32'h3edfbe0c,
32'h3c4000c2,
32'h3e055719,
32'hbf0907d8,
32'h3e121df4,
32'hbe24a073,
32'hbec5815f,
32'hbf2a9635,
32'hbbd1afb5,
32'h3e000ba2,
32'h3d4953f8,
32'h3f3e6df7,
32'h3e773d75,
32'h3dc84e84,
32'h3e84898c,
32'hbd29a8ed,
32'h3d70ea6f,
32'hbe5fbdaa,
32'h3cae0599,
32'hbe27218b,
32'h3dc9cdc8,
32'hbeb5d301,
32'hbea61138,
32'h3dd66cb3,
32'h3e6a3f97,
32'hbea0544e,
32'hbde67207,
32'h3e1a00cf,
32'h3d6cd667,
32'h3dbf9627,
32'h3e3dce88,
32'h3c7f8e13,
32'h3dae967b,
32'h3e9fec11,
32'h3f07e86a,
32'hbee59835,
32'hbeec5ce5,
32'h3e5af521,
32'h3f43b1da,
32'h3e6ee484,
32'hbe333003,
32'h3f12dd41,
32'hbee6cbb7,
32'h3ddf2334,
32'h3e61ad2e,
32'h3e490d18,
32'h3d99bd61,
32'hbc0048c1,
32'h3cdd0f07,
32'hbd90b0a6,
32'h3ed49f98,
32'hbf5abc1a,
32'hbdbc39e2,
32'h3d8b7f31,
32'h3f0dfd0d,
32'h3ec6dd64,
32'h3e4e3517,
32'h3ed64cab,
32'h3d358b24,
32'hbc325f2b,
32'h3f0ff8f3,
32'h3f0423c3,
32'h3db48cb3,
32'hbf39f20b,
32'h3f944459,
32'hbf3ca449,
32'hbf254ef5,
32'h3ed660d6,
32'h3e5181f9,
32'h3ea275b4,
32'hbe98710a,
32'h3f60a4fc,
32'hbb04eff5,
32'hbc5b8c02,
32'hbe5f2f1a,
32'hbc5228f5,
32'h3f0a9527,
32'hbf0dbec6,
32'h3f407d5e,
32'h3d250217,
32'h3f382159,
32'hbec26582,
32'hbd9dd5e2,
32'h3e32682c,
32'h3f51c3bd,
32'h3f903a93,
32'h3ea6f09f,
32'hbeaad073,
32'h3d9967ba,
32'hbca54d0c,
32'h3e91bf2c,
32'h3fc2066e,
32'h3ed73914,
32'hbf03f59a,
32'h3e1ce812,
32'hbf824427,
32'hbf69d849,
32'hbeb68a5d,
32'h3e58b2a3,
32'h3eb5e808,
32'hbf1efa20,
32'h3f03d5c6,
32'h3f02149c,
32'h3ea9f909,
32'h3ee0416c,
32'h3ea112ea,
32'h3e838d49,
32'hbf3ba517,
32'h3f1abb0f,
32'hbdb5cebc,
32'hbe4989a0,
32'hbf855b8d,
32'h3f37a8df,
32'hbf1a5b09,
32'h3ef1c827,
32'h3f1a6012,
32'hbe31fc51,
32'hbe84fcf4,
32'hbdadd007,
32'hbd25de5d,
32'h3d398997,
32'h3ea186fc,
32'h3df1a7b1,
32'hbdb2634c,
32'hbd2d399d,
32'hbf4763bc,
32'hbfa33afb,
32'hbebad1bb,
32'hbf1d716f,
32'h3f7d1814,
32'h3e8f19cd,
32'h3f9dd037,
32'h3daee22a,
32'h3d809d89,
32'h3f42948d,
32'h3f25abc1,
32'h3d96ea6a,
32'hbe9b5260,
32'h3f2777c1,
32'hbec58220,
32'h3f05748e,
32'hbf57882a,
32'h3f476635,
32'hbfdb8882,
32'h3e94bb09,
32'h3f4c458d,
32'h3dc8a403,
32'h3f0d1076,
32'hbd424f75,
32'h3dac2d41,
32'h3ec763ef,
32'h3f3bc983,
32'h3f058f69,
32'h3ea4333a,
32'h3f15c538,
32'hbf0301ee,
32'hbfb1e26d,
32'hbe8edb79,
32'hbeee2f49,
32'h3f4c537f,
32'hbf2516ef,
32'h3fbf537b,
32'h3cbc89e4,
32'hbd8ca825,
32'h3eb168a7,
32'hbe066ed1,
32'h3f5fd9f9,
32'hbd989b4a,
32'h3f349037,
32'hbf09f223,
32'h3f09c96f,
32'hbe90ccd3,
32'hbe9efcc5,
32'hbfb7e8b7,
32'h3f3eb151,
32'h3f1f88a6,
32'hbec780dc,
32'h3ed2fbcf,
32'h3da41a73,
32'hbd322d6b,
32'h3e51c813,
32'h3ea700e6,
32'h3f1836e3,
32'h3e840734,
32'h3e36769b,
32'hbeab7e28,
32'hbfea40f1,
32'h3e70b397,
32'hbf145978,
32'h3f224d73,
32'hbf75e4ad,
32'h3fa221fd,
32'hbf239640,
32'hbf059b1f,
32'h3e642c6b,
32'hbef52f7a,
32'h3f9881be,
32'h3e9051d2,
32'h3e2c293d,
32'hbf3f81b6,
32'h3db82684,
32'hbe0501ff,
32'h3ba0bb82,
32'hbfad43c0,
32'h3f1c7ea5,
32'h3f235619,
32'hbe0fae10,
32'hbeabaa3b,
32'h3be3dc48,
32'h3cc07b64,
32'h3ea21d43,
32'h3eb0cc82,
32'h3f9957f4,
32'h3f41b510,
32'h3e44722f,
32'hbe6039b1,
32'hbff81fd9,
32'h3e1e1b42,
32'h3c94f526,
32'h3f1245af,
32'hbf1df0c9,
32'h3f976efe,
32'hbeb6daa7,
32'hbeb2d1c5,
32'h3f313afd,
32'hbd80c659,
32'h3f514128,
32'h3ea27bdb,
32'hbe91906c,
32'hbe9f2b75,
32'hbf1aed97,
32'hbf233b32,
32'h3eb7964f,
32'h3dcc5af0,
32'h3f86b8db,
32'h3f9a6a1d,
32'hbf155075,
32'h3f62415c,
32'hbdbc6d6e,
32'h3cca3ef1,
32'hbc5d2b29,
32'hbde1a610,
32'h3d92a429,
32'h3ee58e24,
32'h3f229827,
32'hbd71250f,
32'hbf9581f3,
32'h3d936a05,
32'hbf006cea,
32'h3e9c86cd,
32'hbf7ced24,
32'h3f5ef860,
32'hbf0fc273,
32'hbec58459,
32'h3f52844f,
32'h3e1568f9,
32'h3df3a4bf,
32'hbe8a4cd8,
32'hbf5a7d44,
32'hbf026b4b,
32'hbeb1239d,
32'hbf38c6b6,
32'h3e13e927,
32'h3f388b92,
32'h3ebb1e7f,
32'h3f635d1a,
32'hbf70959d,
32'h3f1764fa,
32'h3c737aac,
32'h3d22c306,
32'h3f27d9a1,
32'h3e82503e,
32'h3ed4e9e5,
32'h3e80a5a0,
32'h3f0b4c9a,
32'h3dd352cb,
32'hc040f51f,
32'h3c23dbe5,
32'hbf6fffd7,
32'h3e161f53,
32'hbee5b7b9,
32'h3f2e47e9,
32'hbed2bda6,
32'hbf0211cd,
32'h3e63da5b,
32'hbeb180fd,
32'h3ed9e974,
32'hbee8fc20,
32'hbff4716d,
32'hbf2b6d63,
32'hbf051c1a,
32'h3e1eaa34,
32'h3ee4d760,
32'h3cfdd95e,
32'h3e85b70b,
32'h3f6c1fa6,
32'hbee7dd41,
32'h3d1d8825,
32'h3c7e8ce7,
32'hbd149b1d,
32'h3df9cd87,
32'hbe64e0db,
32'hbe5b00e3,
32'h3eb5b377,
32'h3ee84e04,
32'hbe9519e0,
32'hbf73633a,
32'hbd8c87bf,
32'h3c9bb809,
32'h3e8001d6,
32'hbd2813d8,
32'h3f546cf3,
32'hbe1280b0,
32'h3efefd5f,
32'hbd4eb6d2,
32'hbda697b4,
32'h3f458b67,
32'hbe3fe6d3,
32'hbf925aa9,
32'h3eeae828,
32'hbe342ec6,
32'hbe723ad0,
32'h3ef458ed,
32'h3eca986e,
32'hbeee2bb8,
32'h3f432dbb,
32'hbe9b45ea,
32'h3f4a05c1,
32'hbd957605,
32'hbce8a816,
32'h3b7846bb,
32'hbe031978,
32'hbeb82556,
32'h3ed76a60,
32'h3e9f7674,
32'hbf269c41,
32'hbfb56316,
32'hbd78f3f6,
32'hbf93250c,
32'h3d9208ed,
32'hbe41dc28,
32'h3f3310d0,
32'hbe1c5a44,
32'h3eb0fd00,
32'h3dac777e,
32'h3e30af8a,
32'h3f13840b,
32'hbe80316d,
32'hbead0ea5,
32'h3e81aabe,
32'hbf25777d,
32'h3eb6868b,
32'h3efbdc0a,
32'h3e0c151a,
32'hbf1804bd,
32'h3f51553c,
32'h3ea44971,
32'h3f157dc8,
32'h3d8363ec,
32'h3d721870,
32'h3e40e112,
32'hbdb0f4f1,
32'hbb137866,
32'h3e773a7a,
32'h3e24fb75,
32'hbf09205a,
32'hbf288e7a,
32'h3b4939d9,
32'hbfbcaa77,
32'h3ea921c7,
32'h3ddf6de2,
32'h3f2adfab,
32'h3da5447c,
32'hbe0af679,
32'hbe96c10b,
32'h3f13437c,
32'h3f1963fa,
32'hbe2f8223,
32'h3e064009,
32'hbcbeeb81,
32'hbf2eb614,
32'hbee1e3f1,
32'h3dc0e6bf,
32'h3ebaaaef,
32'h3ed2b21b,
32'h3e569a0e,
32'h3e93ffe6,
32'h3e678f08,
32'hbda45bdc,
32'h3d25d136,
32'h3e5d6c73,
32'h3c6b42a5,
32'h3e94e7b9,
32'h3eca5c8e,
32'h3dca8a8c,
32'hbec45aef,
32'hbdb5371f,
32'hbd9dbbc4,
32'hbecc6edf,
32'h3dd81675,
32'hbd9dc42e,
32'h3f2501ba,
32'h3e8c7f73,
32'hbe9fe705,
32'hbe1548d2,
32'h3ee0ae49,
32'h3f7218e1,
32'hbe31e12b,
32'h3eb4c418,
32'hbdf4f27f,
32'hbf90fa9c,
32'hbf244516,
32'h3d8908b6,
32'h3f3d5893,
32'h3bc52b2d,
32'h3efe481f,
32'hbe0765fc,
32'h3e3676c6,
32'h3db07a04,
32'hbbee021c,
32'hbdc2bf9b,
32'hbcbff91b,
32'h3f075814,
32'h3da5a85e,
32'hbd00376f,
32'hbec6affb,
32'hbeee0f92,
32'hbde6b7da,
32'hbf3ef0fa,
32'h3e8ede99,
32'hbe361058,
32'h3f50abc9,
32'h3ef55c5e,
32'hbe99ed9e,
32'h3d70aca5,
32'h3f2cdd6d,
32'h3ede52f6,
32'hbe600b99,
32'h3e78bf5a,
32'hbdae5f7b,
32'hbecf1ec7,
32'hbf33f4fe,
32'h3ee194ae,
32'h3dd09784,
32'hbe1cdf09,
32'h3e50d6e6,
32'hbde1bf76,
32'hbee172ef,
32'hbd934fce,
32'h3c96b240,
32'hbe0c4d3a,
32'hbea4a9b4,
32'h3f3d796f,
32'hbd431743,
32'h3ed0b51f,
32'h3df8fda7,
32'h3e925489,
32'h3f2f29aa,
32'hbeef381f,
32'h3d874091,
32'h3e105f55,
32'h3f551535,
32'hbed95056,
32'hbe1f8993,
32'hbee323f6,
32'h3efce9d0,
32'hbcc5a178,
32'hbbfbd6f3,
32'h3eca40ba,
32'hbe4b81e6,
32'hbf94865c,
32'hbe5e6398,
32'h3eac2da2,
32'h3b944078,
32'h3eabb093,
32'h3f8e91db,
32'hbeecfe01,
32'hbf1400ab,
32'hbcb05cae,
32'h3db17ff7,
32'hbec78f79,
32'hbeff7634,
32'h3e36bac0,
32'hbdff627a,
32'hbeaab784,
32'hbdb42fda,
32'h3ed07a6c,
32'h3e6a1222,
32'hbee5ebfe,
32'h3ec5198e,
32'h3c5ef219,
32'h3d3b9726,
32'hbebf90d0,
32'h3b8cf080,
32'h3e6a281d,
32'h3f53a344,
32'h3ec48460,
32'hbf2c25ce,
32'h3d9c81ac,
32'hbe3065a3,
32'hbf2b68e5,
32'hbe631e75,
32'h3f574d71,
32'h3e94456a,
32'hbf95a9a2,
32'h3e8866fe,
32'h3d7f231d,
32'hbf469294,
32'hbd10042f,
32'h3ccf1510,
32'h3a9a4e81,
32'hbf2b001f,
32'h3ef4ded2,
32'hbae7c51e,
32'hbef53719,
32'h3ee71980,
32'hbf02c650,
32'h3ecf2ee7,
32'h3f325fc8,
32'h3f232ee1,
32'h3e03d8dd,
32'h3ef7f782,
32'h3d19b84c,
32'hbd519392,
32'h3d31ba0f,
32'h3ebddc92,
32'h3e436ed7,
32'hbf07453c,
32'h3ecabfeb,
32'h3d0760fd,
32'h3d7a8b11,
32'hbf26fe94,
32'h3f423cee,
32'h3da265c7,
32'hbfa5a922,
32'hbe8d8b7e,
32'hbdace00f,
32'h3f8fdcea,
32'hbdd87271,
32'hbc26fe38,
32'hbe888f61,
32'h3f2cb247,
32'hbdba3cc8,
32'h3cf44069,
32'h3f3046d4,
32'h3eeb928c,
32'hbfb3bfba,
32'h3efe744b,
32'hbd1845f2,
32'h3d0ea8c6,
32'h3ec02921,
32'h3eb0cdb9,
32'h3eb558fb,
32'h3e71894f,
32'h3ec5c475,
32'h3c5d7cd7,
32'h3d8d9e3c,
32'hbd85d8d4,
32'h3eacc972,
32'h3ee657f3,
32'h3f72cc76,
32'hbe32acf2,
32'h3f03328a,
32'hbe02ee65,
32'hbfcfbb78,
32'h3f28bebe,
32'h3defe45f,
32'h3c7fa154,
32'h3dd2417e,
32'hbd885b69,
32'hbeb3d0e5,
32'hbf08379d,
32'hbea78ee2,
32'h3e97645d,
32'h3eb9203c,
32'h3e5a1855,
32'hbcf42f8f,
32'hbebbf489,
32'hbe9592e7,
32'hbd5ef0d0,
32'hbf96ba14,
32'h3f75fbf6,
32'hbf133edd,
32'h3c51d19e,
32'h3d3793ee,
32'h3d031e29,
32'h3d4dfde3,
32'h3e6720f4,
32'hbeb4e1cb,
32'h3ebb2758,
32'hbd1043e6,
32'hbe066b40,
32'h3e5cda47,
32'h3eca090e,
32'hbf079ca0,
32'h3ea39974,
32'h3ed8e517,
32'hbd990f91,
32'hbcb12949,
32'hbc0871a3,
32'hbf0929c4,
32'hbde65e45,
32'hbf1a6ebb,
32'h3e6e5582,
32'hbe58d93d,
32'h3edc2c18,
32'h3d5c7769,
32'h3dcc43b6,
32'hbea26b1e,
32'h3f21b5a2,
32'hbf685dbd,
32'h3d30717a,
32'hbe83fc3d,
32'h3d8df95a,
32'h3e873b8e,
32'hbd29bea0,
32'h3e8103e6,
32'hbf00d91b,
32'hbeac8220,
32'h3d8bb51b,
32'hbbd39c67,
32'h3ebbcec1,
32'h3d1947ef,
32'hbebc9cd7,
32'h3e6bc499,
32'h3ebf9fd0,
32'h3f227936,
32'hbdc28f9a,
32'hbd938a2f,
32'h3d49e406,
32'hbd8b04f7,
32'h3f1baad8,
32'h3de34fb5,
32'h3e108cd8,
32'hbddb7751,
32'h3e2165d8,
32'h3dcf28c2,
32'h39e9d550,
32'h3db4f453,
32'hbef13218,
32'hbeb2837e,
32'hbe358f7a,
32'h3db5a56a,
32'h3c6141db,
32'h3d9d914b,
32'hbefdb28c,
32'h3ef9856b,
32'h3e9181a5,
32'hbe30023a,
32'hbd01bbbe,
32'h3dc7b6b9,
32'hbcf1bc24,
32'h3cf7c2e2,
32'hbd788c5e,
32'hbd69dc44,
32'hbdd7067e,
32'h3d0fb3d0,
32'hbd984c27,
32'hbd7ebdf6,
32'hbc18062f,
32'h3e67d443,
32'hbdce07db,
32'hbcaacab4,
32'hbe84ec8e,
32'h3d050351,
32'hbc30f3b4,
32'hbc0813c5,
32'h3d286bf0,
32'hbd983f0c,
32'h3e6b68b8,
32'h3d239363,
32'h3edd1240,
32'hbdbb50dd,
32'h3d1242d2,
32'hbe92d58c,
32'h3c6346a0,
32'hbdccabdc,
32'h3e93c64b,
32'h3d6b5811,
32'hbd57ad57,
32'h3c588091,
32'h3d2c4750,
32'hbd4e3b2b,
32'hbc169125,
32'hbce68f00,
32'hbca74b62,
32'hbd1b5e2b,
32'hbd7d9dda,
32'hbc947d31,
32'h3ae21c70,
32'hbce17117,
32'hbdc13b26,
32'h3c1b705d,
32'h3bc47f11,
32'hbc963135,
32'h3c2050b4,
32'h3cdb97e3,
32'h3dc6a4fb,
32'hbd0e9d33,
32'h3d264ab3,
32'h3d52a016,
32'hbca47d2a,
32'h3d503548,
32'h3bea37d3,
32'hbb2bf99c,
32'h3ce7237d,
32'hbc842a67,
32'hbcef426d,
32'hbdcfc25d,
32'hbc73fd53,
32'hbd8ceeef,
32'h3ccc17e1,
32'hbd32d488,
32'h3d7890f7,
32'hbbd31905,
32'h3d8c501f,
32'h3c613ba3,
32'hbc626bfa,
32'h3d9c7c9d,
32'h3cc24f90,
32'h3d5d148c,
32'hbdd74259,
32'h3d246fe5,
32'hbca13d5b,
32'hbd118f27,
32'hbd04fbe0,
32'hbcacd15d,
32'hbc31fa09,
32'h3d81ec8c,
32'h3d74bc88,
32'hbcfc9ed3,
32'h3ba230e2,
32'h3c0ed4aa,
32'h3d0cb3c8,
32'hbbc3f0ce,
32'h3dca1002,
32'hbd9b1f6f,
32'h3d28a24a,
32'h3d003252,
32'hbb71aeac,
32'h3b888b8b,
32'hbd15d13c,
32'hbd4bef79,
32'h3d418760,
32'hbec3bf1a,
32'hbd3a0f70,
32'h3d7177a0,
32'hbd04325a,
32'h3d199bea,
32'hbd814c09,
32'h3bf1eb89,
32'hbd89a0ab,
32'hbcb3bca6,
32'hbea798d9,
32'hbdb751d6,
32'h3d7baa27,
32'hbbd6b0bf,
32'hbadc6ecc,
32'h3c108f6b,
32'hbe2a4eff,
32'h3cf8e9b2,
32'h3ee44116,
32'hbf0eceb5,
32'h3d8a4c3f,
32'hbf045f3c,
32'hbcb9b459,
32'hbe2905fc,
32'h3e01de07,
32'h3ed88180,
32'h3dc63fc2,
32'h3df649b5,
32'h3d189618,
32'h3d3469f5,
32'h3d8d2d62,
32'h3e50288d,
32'h3e889cb2,
32'h3cdda96a,
32'h3f385336,
32'h3c6c7dd3,
32'hba3e9767,
32'hbe0d02e1,
32'h3e2e05ad,
32'hbd33ac8b,
32'h3f51d7d9,
32'hbcce9aa7,
32'hbc6fa00f,
32'h3c7b2b49,
32'hbc177320,
32'hbe663a05,
32'hbf33ce3d,
32'hbf2d6f0d,
32'hbf828dca,
32'h3d495fc9,
32'h3d4faf2e,
32'h3e4eabda,
32'hbd672299,
32'h3da5b5a3,
32'hbeaf2001,
32'h3ec7e0c8,
32'hbce57bda,
32'hbeaefa94,
32'h3e59cd6e,
32'hbe029652,
32'h3cd499ed,
32'hbe6bf4bb,
32'h3f48a42c,
32'hbd9e12ef,
32'h3f38123d,
32'hbd6fc929,
32'hbd2b7886,
32'h3c88ad4e,
32'hbeac2754,
32'h3e12e28e,
32'h3f26a534,
32'hbd87d3df,
32'hbf09b162,
32'h3e83dffc,
32'hbe8f05a3,
32'hbdab5b01,
32'h3f209573,
32'hbf293092,
32'h3ad80450,
32'hbf04566e,
32'h3e9fd5f1,
32'h3e086b05,
32'h3e9fcd0c,
32'h3e199e1b,
32'hbf80f0b2,
32'hbe88a266,
32'hbead0c38,
32'h3e386b38,
32'h3ec6dce3,
32'h3f10bbc3,
32'hbeba4e8d,
32'h3f499665,
32'h3e3d04ea,
32'h3e9fadb4,
32'hbcdea8bc,
32'h3bb3c810,
32'hbc9325eb,
32'hbf9fa39d,
32'h3e4895dd,
32'h3f17ecfb,
32'hbe8f9c42,
32'h3ec77164,
32'hbe3277a7,
32'hbf0fb15f,
32'h3e1f23fb,
32'h3e1d5912,
32'h3edb6b57,
32'h3c88fe77,
32'h3f1b488f,
32'hbdb02c54,
32'h3e127620,
32'h3f22ec14,
32'h3f39eaca,
32'h3e94fb55,
32'h3df40726,
32'hbe836096,
32'h3dec5406,
32'h3dc8366d,
32'hbf28d19d,
32'h3f0fb496,
32'hbf19d854,
32'h3fa8bc3f,
32'h3e9eb817,
32'h3dfd2d0c,
32'h3f32c845,
32'hbc515cc7,
32'h3d1010de,
32'hbf8903d7,
32'hbefb40bc,
32'h3f33cdb0,
32'h3e1c31e0,
32'h3f160e18,
32'h3f3d7a33,
32'hbcb3c3b4,
32'h3f434ab0,
32'h3f135cbd,
32'hbe7c7985,
32'hbe559f57,
32'hbf409670,
32'h3f62b598,
32'h3f1d0cc3,
32'h3efe0bf6,
32'h3f564793,
32'h3dcc34c2,
32'hbe8a89f2,
32'hbe411094,
32'h3ec69f44,
32'h3eb884e8,
32'hbf336ca4,
32'h3f03b8bf,
32'hbf88c270,
32'h3f359c52,
32'h3ea587ad,
32'h3f1f62e0,
32'hbe3647fc,
32'h3b8de391,
32'hbc0f6a61,
32'h3d71825f,
32'h3e611199,
32'h3eb04012,
32'hbf09b262,
32'hbc995252,
32'h3e68e7be,
32'h3d80ee9a,
32'h3e326e06,
32'h3e85801d,
32'h3e744abe,
32'hbee499e8,
32'hbe888c98,
32'h3f0c4877,
32'h3f3decd7,
32'h3d623b7c,
32'h3f34eafb,
32'h3cadec3f,
32'hbf88fb10,
32'h3f3a6a9e,
32'hbf93d6d6,
32'h3f20618e,
32'hbee8663c,
32'h3f237a26,
32'hbfab021a,
32'h3cae4719,
32'hbe0bf939,
32'h3e684e4c,
32'h3f1804a8,
32'h3d09d079,
32'hbd54c4a3,
32'h3dbc4588,
32'h3f06a258,
32'h3ea3b197,
32'hbca7b001,
32'h3f3bef27,
32'h3f56a1a2,
32'hbdd319bf,
32'h3e393d6a,
32'h3f0fa5d5,
32'h3f003adc,
32'hbfb87230,
32'hbea87179,
32'h3f135883,
32'hbf075775,
32'hbcc5c547,
32'h3eb4493b,
32'hbe5ef861,
32'hbf25266c,
32'h3eedc9cc,
32'h3e81ec97,
32'h3ee5b650,
32'hbe32c0ff,
32'h3f7126af,
32'hbf6107cf,
32'h3f694a0f,
32'h3d709145,
32'h3f239151,
32'hbe269214,
32'hbd86f83c,
32'h3aa65781,
32'h3ea8daaf,
32'h3dd59a99,
32'hbeee76e1,
32'h3ea450fd,
32'h3e45d651,
32'hbe8a2d70,
32'hbeea50b2,
32'h3d903fa9,
32'hbe65f054,
32'h3ea5e60f,
32'hbeb1721f,
32'h3ed73d75,
32'h3eb1eaf5,
32'hbe2f0d6b,
32'h3d831772,
32'h3eb446f0,
32'h3e617b88,
32'hbf12e51e,
32'h3eaf9ce2,
32'hbdab9276,
32'h3e258f8f,
32'hbebc2d53,
32'h3e899487,
32'hbc58a35e,
32'h3e789fe8,
32'h3e150232,
32'hbe899f8a,
32'hbf28a645,
32'h3d34df63,
32'h3d2ed010,
32'h3eb1ceda,
32'h3ecc08b8,
32'hbe24bb8f,
32'h3ec270ee,
32'h3e0f3c2f,
32'hbe92e510,
32'hbf981c73,
32'hbc605a4d,
32'hbeabf692,
32'h3ebc4201,
32'h3ca9570f,
32'h3f020878,
32'h3ecc6123,
32'hbf40512e,
32'h3d5ba9e5,
32'h3e63ba3c,
32'h3edfdeb2,
32'hbe01e961,
32'hbefa4a0d,
32'hbf091085,
32'hbe86f288,
32'hbe8899a6,
32'hbf7a50d5,
32'h3ed2834a,
32'h3f0044e0,
32'h3ebb9b1e,
32'hbe2ddaab,
32'h3e4a8239,
32'hbd94abc0,
32'h3d15972b,
32'h3f03df5d,
32'h3ee98218,
32'hbe8ef961,
32'h3df60fac,
32'h3d12755c,
32'hbd980080,
32'hbf3a374e,
32'h3de24bc8,
32'hbf189ac7,
32'h3dc93647,
32'hbf0edd3d,
32'h3d9431c5,
32'h3e3d35c0,
32'hbf1dc298,
32'h3e881bc2,
32'hbe295ebe,
32'h3e68c7ef,
32'hbe82fd28,
32'hbecdc9fc,
32'hbebada00,
32'hbeceec8f,
32'h3dee7904,
32'hbf606186,
32'h3ecd398b,
32'h3ef695e3,
32'h3e3beaec,
32'h3eb6f5e6,
32'h3eb0bdf0,
32'h3b5a60b8,
32'h3d893e18,
32'h3ea87551,
32'h3e9d8eae,
32'hbe7def7c,
32'h3e1ce811,
32'h3f0d3e78,
32'h3e69c9f0,
32'hbe8295ae,
32'h3e86a56d,
32'hbf125c80,
32'h3e182c82,
32'hbf44ac53,
32'hbe13444e,
32'h3eb9468b,
32'h3e1cc642,
32'h3eba5f4a,
32'hbeaf9143,
32'h3ede2a93,
32'hbf1c3c2f,
32'hbea7bdfb,
32'hbe701c3f,
32'hbda72345,
32'hbe2fb6e7,
32'hbf3fd0a3,
32'hbe150aa3,
32'h3edc5cf7,
32'h3e36ebcf,
32'hbe3de130,
32'h3cf8c206,
32'h3d3e2da8,
32'hbce7b1b7,
32'h3c20387b,
32'h3f20b09b,
32'hbe58d355,
32'h3e94a23e,
32'h3f07aaf8,
32'h3e2dc489,
32'hbcbd6888,
32'h3ee2165c,
32'hbf093da0,
32'h3e33eada,
32'hbeea9bc2,
32'hbb5acc34,
32'h3ce4ebd3,
32'hbe418eb8,
32'h3e6f8823,
32'hbeffcbc9,
32'h3e1a6a86,
32'hbf0c5cfe,
32'hbf79b7e9,
32'hbe5ba880,
32'h3ec72aa3,
32'h3e143f92,
32'hbe8c87df,
32'hbe0628c4,
32'h3e214690,
32'h3e49b9f9,
32'hbf78b1f0,
32'h3de60492,
32'hbca8fc00,
32'hbd111d51,
32'h3d939406,
32'h3e42a9e6,
32'hbe99844a,
32'h3e685c2f,
32'hbd2132d2,
32'h3e216cd2,
32'hbf145d15,
32'hbd470d7d,
32'h3d2ff62b,
32'hbd3cd1b1,
32'hbefcbd24,
32'hbdd12051,
32'hbe9c5c89,
32'hbeec661e,
32'h3df46677,
32'hbe4a8fe6,
32'h3debd9b6,
32'hbebc542c,
32'h3d5ee7fd,
32'hbea5acf8,
32'h3e324a4e,
32'h3b92d7c1,
32'h3d35a2e5,
32'h3d833e50,
32'hbc0e485f,
32'h3e41349d,
32'hbf7aeffb,
32'h3c3bab35,
32'h3d5b7f70,
32'h3db9f7f4,
32'h3e43c341,
32'h3e38ac9b,
32'hbdf0768e,
32'h3e19bee9,
32'h3dac4d3c,
32'hbf357149,
32'hbfb8d8e0,
32'h3e9e9140,
32'hbb62c9d2,
32'h3da64605,
32'hbe87289b,
32'hbe0b940b,
32'hbe484936,
32'h3ee8703a,
32'h3e9a1f87,
32'hbe53a1f5,
32'h3e6aaaa3,
32'hbed69381,
32'h3f5d653a,
32'hbf1004f3,
32'hbd00b8f5,
32'h3d04152e,
32'hbefd9a5b,
32'h3dd55dea,
32'h3da7b2bb,
32'h3e497450,
32'hbf22f8ac,
32'h3e114c6b,
32'hbe1b44ce,
32'h3c85f6e1,
32'hbde6e79c,
32'h3b861905,
32'h3ded9c38,
32'h3e06aef2,
32'hbea22dc4,
32'hbf7e38b8,
32'hbf8cb9e4,
32'hbeb2ebe2,
32'hbf1cea35,
32'h3e4deb74,
32'hbe089f1b,
32'hbe3321fd,
32'h3d92c249,
32'hbe355f14,
32'h3e2d5fc4,
32'hbe790e2b,
32'h3e9adcb9,
32'hbe36a975,
32'h3e88d360,
32'hbd073a33,
32'hbe4898ae,
32'h3e6e0468,
32'hbf3cc0f6,
32'h3c0ce3bc,
32'h3e105cb7,
32'hbc1af71a,
32'h3d8c238d,
32'hbe23ec4e,
32'h3c9c7069,
32'hbd8ebf3b,
32'hbea9473e,
32'hbd6542d3,
32'h3e050385,
32'h3e210acb,
32'h3e90aaf9,
32'h3cf928bf,
32'h3c29ef33,
32'hbecad1c2,
32'hbcebf2de,
32'h3e7a9d4c,
32'hbe20cc36,
32'hbdd0bbbf,
32'hbe004436,
32'hbeaf9777,
32'h3d9e0910,
32'hbdd9879d,
32'h3edbb6e3,
32'h3e38edca,
32'h3e1fe441,
32'hbe4c9832,
32'hbe7f2b02,
32'hbd8eac25,
32'hbf4f8479,
32'hbd628878,
32'h3e242771,
32'hbe849b5d,
32'h3e8f9196,
32'h3e52e7f0,
32'hbda446ea,
32'h3bd2e170,
32'hbe74b298,
32'h3e870441,
32'hbe0c7604,
32'h3dc59a92,
32'hbd0009ea,
32'hbefae1e3,
32'hbeeb4b28,
32'hbda97cd5,
32'h3cbf889e,
32'h3e89d4b4,
32'h3e4dbb41,
32'h3e0f47d5,
32'h3d279b64,
32'h3d80eb42,
32'h3e127f42,
32'h3e2fc8f1,
32'h3f08d80e,
32'hbe8648df,
32'h3e5ae81b,
32'hbeb38b01,
32'hbdfa207e,
32'h3eeba15f,
32'hbe75b0b9,
32'h3ec8436f,
32'h3dd1701d,
32'hbd61c901,
32'hbdbaa92b,
32'h3dd84173,
32'hbcc49524,
32'hbdd0d8b5,
32'h3c54b93c,
32'h3e94db20,
32'h3d876fd4,
32'hbe9af8cd,
32'hbe0c20f3,
32'hbe660ff8,
32'hbebc6071,
32'hbef959ae,
32'hbecc7778,
32'hbb56782a,
32'hbed881f8,
32'hbd413ad0,
32'h3d9162e0,
32'hbf8356fc,
32'h3b7bce35,
32'hbde72737,
32'h3e9559d7,
32'hbbfc2182,
32'h3f0cf4a3,
32'h3eb3a1c3,
32'hbea36c3c,
32'h3d70e93f,
32'h3eb7d9ad,
32'h3d294451,
32'hbe3c73c5,
32'hbe286fde,
32'hbe30492e,
32'hbf027bad,
32'hbc138101,
32'h3c941642,
32'hbed3c67d,
32'h3e361d9e,
32'hbdeeb77a,
32'h3cc1a858,
32'h3ee2b92a,
32'hbdba89e7,
32'h3eef59cb,
32'hbd48f6e2,
32'h3ed9c29d,
32'hbe9354f4,
32'h3e50ca3e,
32'hbe7f25a6,
32'hbd992a61,
32'hbe5256ca,
32'h3cf4b7f6,
32'hbe8d8bc3,
32'h3d5e5f84,
32'h3d92d1eb,
32'h3f33c96c,
32'h3d31ffd8,
32'h3e90c863,
32'hbe4d701c,
32'h3f2aaac1,
32'hbe6e06f9,
32'hbec4e92b,
32'hbc9818da,
32'hbe981f62,
32'hbf4014ec,
32'h3dac2a68,
32'hbcce57dc,
32'hbed96570,
32'hbd78b012,
32'h3dcc0a3a,
32'h3e0e7683,
32'h3de10a0e,
32'hbda32059,
32'h3e8df6c0,
32'h3e635e88,
32'h3e2f2ac9,
32'hbc1c26f5,
32'h3edf888b,
32'hbd3eb8b3,
32'h3d0b2ba4,
32'hbedb5988,
32'h3e2654ab,
32'hbe14c737,
32'h3d08f1e1,
32'h3e1e5cf0,
32'hbdc9ad68,
32'h3deeff85,
32'hbe441e4b,
32'h3d9a5411,
32'h3f863b4d,
32'h3e5fee2b,
32'hbf014428,
32'h3d3e9538,
32'hbee74ac0,
32'hbf296707,
32'hbd96b34b,
32'hbd1cf16e,
32'hbb891d28,
32'hbeabeb58,
32'hbe49bd41,
32'h3c3e3e56,
32'hbf293750,
32'h3f19fad4,
32'h3e75721d,
32'h3ec78413,
32'h3ea3998f,
32'h3f080b3f,
32'hbdedd3e0,
32'h3e28ed84,
32'hbecef980,
32'hbebced8a,
32'h3ec7949c,
32'h3da8372a,
32'hbd27468a,
32'h3ef36806,
32'h3ee4921d,
32'hbe2ffec1,
32'hbe2543ea,
32'h3e1b53f5,
32'h3f9e3959,
32'h3ec2d538,
32'hbece388b,
32'hbdcc45aa,
32'hbefe4574,
32'hbebf2cf9,
32'hbd15ecb0,
32'h3cacc572,
32'hbd771582,
32'h3eab76ec,
32'h3e8c90d4,
32'hbe3f261d,
32'hbe2f11f7,
32'h3f60de3d,
32'hbc707b42,
32'h3f52dc3c,
32'hbed1f335,
32'h3db33f0c,
32'h3de97ade,
32'h3e5a7250,
32'h3f039f39,
32'hbeed1a79,
32'h3efa94a0,
32'h3e19fa00,
32'hbeba4c22,
32'h3e78b8cc,
32'h3cb81c2c,
32'h3e35a404,
32'h3f161d88,
32'hbe2d6f07,
32'h3f5c9f2d,
32'h3f0f579a,
32'hbec2afd2,
32'hbe83e17a,
32'hbed8390e,
32'hbf12d9e6,
32'h3b34e5d1,
32'h3ccf6256,
32'h3d88b939,
32'hbf346714,
32'hbf0acca3,
32'hbe710ad6,
32'hbea43102,
32'hbe4ad751,
32'h3e7ff6bd,
32'h3f2443de,
32'h3f266082,
32'h3ec1a9a3,
32'hbe0635cd,
32'h3eb24258,
32'hbf6cdcae,
32'h3d874090,
32'h3f2109d5,
32'h3eb933ce,
32'hbe867027,
32'h3e12a87b,
32'hbf15d23c,
32'h3ee10751,
32'hbeb9c4c7,
32'hbe53f70c,
32'hbd11175f,
32'h3ea274c1,
32'hbeaa933f,
32'hbd57341a,
32'hbed1f0f6,
32'hbe3596b6,
32'hbd0a0cb8,
32'h3c22b9b0,
32'hbe373205,
32'hbfabd716,
32'hbfbda1a9,
32'hbf31ac9b,
32'hbf2a8f48,
32'hbe8c40ad,
32'hbe99b3e9,
32'h3eadd15e,
32'h3ed5acbb,
32'h3f753899,
32'hbfc18f19,
32'h3eab7324,
32'hbedffa30,
32'hbd46cf76,
32'h3f7285f6,
32'h3ee27030,
32'hbefe3a35,
32'hbe9f1a77,
32'hbf65b36d,
32'h3f083025,
32'hbf469fad,
32'hbf04371f,
32'h3f905311,
32'h3ed62d1a,
32'h3eea1975,
32'hbebbe44f,
32'h3f4515f0,
32'hbbdcfdde,
32'hbcb1de19,
32'hbdd5feca,
32'h3e394e98,
32'h3e52f71b,
32'hbf81e3b7,
32'hbed44fa5,
32'hbf93a0c9,
32'h3f09ffe1,
32'h3f812004,
32'h3f8d284b,
32'h3e3e0808,
32'h3ef49bb7,
32'hbed91f88,
32'hbed3c532,
32'hbd417f02,
32'hbd565e8a,
32'h3f2ced5b,
32'h3f0cdf26,
32'h3ea4178f,
32'hbf7a0719,
32'hbe7523fd,
32'h3c657365,
32'hbe3f33e5,
32'hbe9ffe78,
32'h3f077bb7,
32'h3f36ba93,
32'hbb36d617,
32'hbede004a,
32'hbcdf69ef,
32'h3d2ddeda,
32'h3d101576,
32'hbd2db8ce,
32'h3ea068be,
32'hbd82a2f2,
32'hbe019404,
32'hbcfdb00f,
32'hbf057aa6,
32'h3e50d86f,
32'h3d310090,
32'hbc199679,
32'hbe7ce5c1,
32'h3ea316b1,
32'h3d74d5fd,
32'hbed6b702,
32'hbd0db376,
32'h3c990b1c,
32'h3f4f9161,
32'hbefecdd8,
32'hbdd57f5e,
32'hbf4873ac,
32'hbd4cc625,
32'hbda259f0,
32'hbe567c55,
32'hbd44eaa2,
32'hbd8c2710,
32'h3e7a27ac,
32'hbcd2f216,
32'hbd8ed63d,
32'h3d9997d7,
32'hbd7f43f1,
32'h3cf9a9d0,
32'h3ca2938d,
32'h3f388605,
32'hbe3d889c,
32'hbe041e27,
32'hbebd1250,
32'hbee46eeb,
32'hbe3473b3,
32'hbd04f827,
32'hbd8e7562,
32'hbe91119f,
32'hbcb403aa,
32'h3d6868ad,
32'h3e9a4838,
32'hbd562071,
32'h3d745215,
32'hbe23b0f3,
32'hbd9af209,
32'hbd0c7e63,
32'hbdd7d4af,
32'h3dc84925,
32'hbda7af1a,
32'hbd8f6a18,
32'h3cdc9ae0,
32'hbd506140,
32'hbd861a90,
32'h3c9ce572,
32'h3d9d9cd5,
32'hbd85bfc3,
32'h3d24c129,
32'h3c0ca800,
32'h3d2c5c2a,
32'hbd471ee2,
32'hbdaa5c82,
32'h3d84c1d4,
32'h3bbf6c74,
32'hbc9a2e62,
32'h3d52b0bd,
32'hbbba52ae,
32'h3b8274e6,
32'h3d9084b6,
32'hbd461eea,
32'h3b055c6b,
32'hbd5c0583,
32'h3d8e4c6f,
32'hbd87577f,
32'hbd292aaa,
32'hbda73a60,
32'h3d29e4cc,
32'hbcd61907,
32'hba98386c,
32'hbb98e2fa,
32'h3d237dae,
32'h3da45938,
32'h3c4861e5,
32'h3dd0fcbd,
32'hbd754c95,
32'h3d602369,
32'hbdd30219,
32'hbd5b840b,
32'h3de0798b,
32'hbad7007c,
32'hbc3928ff,
32'hbd74826c,
32'h3d0aaf43,
32'h3dbd1fc6,
32'h3da26ab8,
32'hbc9c6f4a,
32'h3d617031,
32'hbdb5ce45,
32'h3c9cf35d,
32'hbd9b2211,
32'h3db37e03,
32'hbdde84b5,
32'hbd1980d7,
32'h3d9c6657,
32'hbcc00ff5,
32'h3cd1291a,
32'hbd301846,
32'hbd0827ee,
32'h3ee2953d,
32'hbde1421f,
32'h3ef51272,
32'hbe29c144,
32'h3c902c2e,
32'h3cca9e38,
32'h3e90cd26,
32'h3e83864c,
32'hbdc08b85,
32'h3f4ff8e5,
32'h3ce9c427,
32'hbd178243,
32'hbe939738,
32'h3f468c90,
32'h3ed73666,
32'h3f696519,
32'h3e39776f,
32'hbdbe05c0,
32'h3c8172c3,
32'h3cb8835e,
32'hbe8af1b7,
32'hbe0455e3,
32'hbf38d9b1,
32'hbf7b8f91,
32'h3eddd945,
32'hbd50399a,
32'h3e5e49bd,
32'hbd7b50c6,
32'hbc18595e,
32'hbed96433,
32'h3f4a96b3,
32'hbe58102a,
32'hbe9e2a20,
32'h3e5bf666,
32'h3e629dd6,
32'h3cc4035d,
32'h3f16309f,
32'h3e751036,
32'hbe791dd9,
32'h3f1aae7a,
32'h3ca12025,
32'h3d9e422e,
32'h3e2ceec0,
32'h3e10d84d,
32'h3d9b0c93,
32'hbd8e6fee,
32'h3e99b559,
32'h3cee8d41,
32'h3e6d7599,
32'h3bf56539,
32'hbe55c054,
32'h3c62527c,
32'hbf1db886,
32'hbe6f7319,
32'h3f6c4551,
32'h3f17397e,
32'h3f7467d1,
32'h3e02f0d7,
32'hbe7d474d,
32'hbf5f07ba,
32'hbd8fe5bc,
32'hbecca205,
32'h3f22f189,
32'h3f4c3e6c,
32'h3ed4c942,
32'hbf04fda1,
32'h3f842356,
32'h3edcee04,
32'h3d405752,
32'hbf5bf1d8,
32'hbdb9f79e,
32'hbbbdd3f7,
32'hbf62b3a4,
32'h3f0d6cf4,
32'h3ee7c059,
32'hbef78d26,
32'h3ec32e77,
32'h3e062da4,
32'hbfba26c4,
32'h3e1f9248,
32'hbd2e72eb,
32'h3e6ed209,
32'hbdbfb5bd,
32'h3ef10ccd,
32'hbd10f13c,
32'hbec6f796,
32'h3dea57ab,
32'h3f2f53bf,
32'h3bb40fda,
32'hbc67127d,
32'h3e911a76,
32'hbf141d46,
32'hbf8cb376,
32'hbf4564ba,
32'h3daddd10,
32'hbfab6e47,
32'h3f5a8be8,
32'hbed2b23e,
32'hbe5f176f,
32'h3e7d09ce,
32'h3d700a73,
32'hbd587812,
32'hbf08dcbf,
32'hbf047f07,
32'h3e947456,
32'h3e5220c6,
32'hbed01e01,
32'h3e14c7cd,
32'hbf10ae68,
32'h3d96b508,
32'hbea72de1,
32'h3e802a5e,
32'hbf248fc8,
32'h3e58de7a,
32'hbea25ef1,
32'h3d8300a9,
32'hbea7ca98,
32'h3ecb6536,
32'hbe956391,
32'hbe6877a0,
32'hbe8bc00d,
32'hbfbe54c6,
32'hbf184bbe,
32'hbe33c962,
32'h3e8a84d9,
32'hbf8c2e2b,
32'h3f04f761,
32'h3d31966a,
32'h3eb766fb,
32'h3ea4cdef,
32'hba9378fa,
32'hbd0a8d2f,
32'h3eb61947,
32'h3e98b252,
32'h3db6201b,
32'hbda33e0e,
32'hbe2bfa97,
32'h3dc41a2c,
32'hbf81c8c3,
32'h3e25c05e,
32'h3d7dece7,
32'h3edcaecf,
32'hbf8bfc16,
32'h3e2870a3,
32'hbec98eb3,
32'hbf178b49,
32'hbf19d0ca,
32'h3e38a3a7,
32'h3d871e3d,
32'hbf587907,
32'hbe53e197,
32'hbfb9b4e7,
32'h3ed04516,
32'hbe6e1c4e,
32'h3f3d2f52,
32'hbe1c44c0,
32'h3e5df566,
32'h3e1ccf02,
32'h3e891d76,
32'hbe145d45,
32'h3a2814ec,
32'h3dae6d7b,
32'h3cf1ea14,
32'h3e8b6fa3,
32'hbe978f23,
32'hbe92e884,
32'h3ec93e1d,
32'h3cc81c7f,
32'h3dc6ae7e,
32'hbcea3516,
32'h3ef4af77,
32'h3e6b8e85,
32'hbfbe3940,
32'h3f086f44,
32'hbd9e8462,
32'h3d5518b4,
32'hbf22ef9c,
32'hbdf88a74,
32'hbe38297c,
32'hbf3dd70c,
32'hbfc459df,
32'hbdcd63bf,
32'h3e4cf8c9,
32'hbe4bcf60,
32'h3f868eb4,
32'hbc674040,
32'h3cb25e47,
32'h3db94f11,
32'hbe035260,
32'hbf46ea09,
32'h3d716cbf,
32'hbd6c35ef,
32'hbd272f4e,
32'hbc5894bf,
32'hbeda164b,
32'hbdfad68c,
32'h3d9cbf95,
32'hbef2c79e,
32'h3f0b45f2,
32'hbe7abfad,
32'h3e5feb84,
32'h3ef4f995,
32'h3f34ed8e,
32'h3e34c784,
32'hbe3f071a,
32'h3f51f566,
32'hbe2a5f0f,
32'h3d0f32a0,
32'hbe857433,
32'hbf00a7fe,
32'h3db5ebf6,
32'hbdaa13d8,
32'h3e8966b2,
32'hbe645b43,
32'h3f3a2c31,
32'hbe4c66d8,
32'hbde269ed,
32'h3ecb7d98,
32'hbeafa959,
32'hbf153495,
32'hbd56c0fc,
32'h3d952ec2,
32'h3df1e14f,
32'h3e77d5ea,
32'hbf21c742,
32'hbdfd9fd1,
32'h3e13b151,
32'hbdd23c07,
32'hbeb3dd53,
32'h3dc3a150,
32'hbe81fed1,
32'h3e817849,
32'h3e81dcea,
32'h3e6860de,
32'hbe900f12,
32'h3ef207a7,
32'h3ca4e41e,
32'hbef33e74,
32'h3db916d2,
32'hbec01a91,
32'hbfd987ab,
32'hbfa1398d,
32'h3e35ed34,
32'hbe3c4c22,
32'h3ea3f24b,
32'h3ee7ecf1,
32'h3d1039af,
32'h3e47476d,
32'hbe2e54e8,
32'hbef4f2f8,
32'hbd903819,
32'hbd3e41a4,
32'h3eb9f0de,
32'h3e63d5ae,
32'hbe912d78,
32'hbda783e6,
32'hbec3ebc3,
32'h3e5c224d,
32'hbe8ca656,
32'h3c94437d,
32'hbe25b539,
32'hbd5d71ed,
32'hbdf3096c,
32'hbe8b674e,
32'hbe91a3c8,
32'hbeb4b51d,
32'hbe64973c,
32'hbcac4985,
32'h3e240004,
32'hbe3ea7dc,
32'hbfd899c1,
32'hbe6c19c6,
32'hbc83be6f,
32'hbe46ed95,
32'hbe301679,
32'h3d8728b3,
32'h3dd2f21f,
32'h3d80b3fb,
32'h3e806c0d,
32'hbd8cf343,
32'hbcc1b339,
32'h3cfcd1af,
32'hbe58d396,
32'h3e0ca114,
32'hbea541ed,
32'h3db65696,
32'h3db76bc5,
32'hbc710e08,
32'hbd119c40,
32'hbdad0b72,
32'hbd6b4e7f,
32'h3d9f7087,
32'hbe4c2fb7,
32'hbd99178f,
32'h3d8655f6,
32'hbe633148,
32'h3e3cf3cf,
32'hbdaaba1b,
32'h3e510ea1,
32'hbebdfee6,
32'hbf6d6871,
32'h3c347933,
32'h3e7b8c4b,
32'hbcd37da1,
32'h3dfec403,
32'hbd43e353,
32'h3dc538c8,
32'h3ee86241,
32'h3e5db391,
32'hbdadf3eb,
32'h3c80e3de,
32'hbd0f8dd1,
32'h3d993245,
32'h3e5ba4b4,
32'hbe7c5956,
32'hbdd3520d,
32'h3e8c3c8a,
32'hbc917b17,
32'h3e3f84cf,
32'hbe9e49d2,
32'h3d3dc34e,
32'hbccb6a35,
32'hbdafff95,
32'h3def5927,
32'hbe534e99,
32'h3df2b923,
32'hbda548b2,
32'hbe217e3d,
32'h3d1a9303,
32'hbf450cbe,
32'hbf808ceb,
32'hbf10cd7b,
32'h3df4074a,
32'hbd51512d,
32'hbdc109d4,
32'hbdabae92,
32'h3e665ec3,
32'h3ea2ddd5,
32'hbb9c1292,
32'hbe6cdd72,
32'h3d77c834,
32'hbdb3f47b,
32'h3e6c7641,
32'h3eaec459,
32'hbe171e6a,
32'hbde2b44e,
32'h3e603181,
32'hbdecf52f,
32'hbeb3eb97,
32'hbea34aeb,
32'h3e30e48a,
32'hbe15bdc2,
32'hbe92de2d,
32'h3e359bd7,
32'h3c3028e9,
32'hbedc41f1,
32'hbe7d0166,
32'hbe08f099,
32'h3d4ff6b2,
32'hbec78978,
32'hbed88d35,
32'hbe99924a,
32'hbe3b8128,
32'h3cce901f,
32'hbd2348c2,
32'hba8d8c76,
32'hbd87dd5a,
32'h3dc7918c,
32'hbec9b186,
32'hbd8b07ee,
32'hbdca8b7f,
32'h3c9815de,
32'hbe2a2ff2,
32'h3e99c744,
32'hbeaaf182,
32'h3d5010e0,
32'hbdbc1455,
32'hbf90155c,
32'hbe813648,
32'h3dff1ec8,
32'hbd24b4fe,
32'hbcd55cc7,
32'hbe781ef8,
32'h3daa9fa8,
32'hbda88a9f,
32'hbee83e89,
32'hbcf1affc,
32'hbced0132,
32'h3e9892bf,
32'h3e6e5426,
32'h3e8b3646,
32'hbf6e9b30,
32'hbd85694c,
32'h3d8893af,
32'hbe402689,
32'hbd819004,
32'h3e35d238,
32'h3e8a4e41,
32'hbe9f3b56,
32'h3e7671b1,
32'hbe19966f,
32'hbb84d55c,
32'hbf000e33,
32'h3e79954e,
32'hbeac9ebf,
32'hbcf6b99a,
32'hbed5fe6b,
32'hbf5526e5,
32'hbd7247f7,
32'hbe724de6,
32'hbeaa24d8,
32'hbd76106a,
32'hbe9fa8fd,
32'h3c3629f2,
32'hbd8e1446,
32'hbe8bf07e,
32'hbeb16445,
32'hbf04247c,
32'h3e099594,
32'h3e60ea52,
32'hbdfc5013,
32'hbf2e30f5,
32'h3e056708,
32'h3e2eea98,
32'hbf079be1,
32'hbb9e933e,
32'hbd535270,
32'h3e8269f7,
32'hbcfa491e,
32'h3e6c4c65,
32'h3d3d71e0,
32'hbb06d4c2,
32'hbf004b1d,
32'h3e9b318f,
32'h3e36db33,
32'hbdbc3112,
32'hbe7b4ab5,
32'h3e88cd91,
32'hbe34eb46,
32'hbdaaa994,
32'h3ec87aa5,
32'h3e312451,
32'hbf0e4b52,
32'h3d5fcd65,
32'hbe2b470a,
32'hbf28c0f5,
32'h3e0b7494,
32'hbe370247,
32'h3e2d7f68,
32'hbead3f16,
32'hbdfc206b,
32'hbf8c23f0,
32'hbe2dd185,
32'h3d176952,
32'hbf26d526,
32'h3e26a623,
32'hbe06b52c,
32'hbe491e7a,
32'hbe2928a2,
32'hbda2ab90,
32'h3ba06421,
32'h3b615e60,
32'h3d8c5c43,
32'h3d528f10,
32'h3e0c1f3b,
32'hbe287c91,
32'hbe836ffa,
32'h3ec97596,
32'hbf23fe88,
32'h3e7cb7a5,
32'h3eadc390,
32'h3e7c844b,
32'hbd78b59b,
32'hbc847689,
32'hbd9dfcce,
32'hbf145cec,
32'h3e7b748b,
32'hbe62e77a,
32'hbdc2b9eb,
32'hbd877ad6,
32'h3c775804,
32'hbfc7123b,
32'hbe46023b,
32'h3c232c44,
32'hbebb2c3a,
32'h3d987ef4,
32'hbc6bc8e4,
32'h3e17f0cc,
32'h3e13886d,
32'hbed703f3,
32'hbd3df73b,
32'hbce18bfb,
32'hbdc1052f,
32'h3d08a4f3,
32'h3e397345,
32'hbd526588,
32'h3e82dbbc,
32'h3e08896f,
32'hbe8ed740,
32'h3e9f863e,
32'hbf06044a,
32'hbe6fc71a,
32'hbbc9f5df,
32'hbdf06a6d,
32'hbdf122ce,
32'hbf4c9160,
32'h3e6ac0a9,
32'hbf014c4e,
32'h3d9c6110,
32'h3e2a896e,
32'h3e248de9,
32'hbf904243,
32'hbe3c48e0,
32'h3e9ab2b4,
32'hbdbff239,
32'h3e38df0d,
32'hbcb60d6f,
32'h3e3b68af,
32'h3edf7286,
32'hbec4b0dd,
32'hbd6cdef3,
32'h3d8514e4,
32'h3b9c0876,
32'h3ea0e282,
32'h3e8972eb,
32'hbe3d5b20,
32'h3d1f3fbd,
32'h3e33655b,
32'hbd60d031,
32'h3ed37ac3,
32'hbea1cc51,
32'hbea977e3,
32'h3c3f735d,
32'hbd04b5ac,
32'hbeb1036a,
32'hbfede605,
32'h3e4a8f47,
32'hbf2ecce5,
32'h3edb9e38,
32'h3e76c90d,
32'hbcab931e,
32'hbf7b4681,
32'hbe6c744a,
32'h3bbff371,
32'hbda88fee,
32'h3e11d173,
32'h3cee8fda,
32'hbdd8fe8a,
32'h3eac8e39,
32'hbfd9c407,
32'hbd4f5cae,
32'hbdd7a028,
32'hbdaed6b9,
32'h3e3e9b59,
32'h3e9ec0c4,
32'hbe4a2192,
32'h3ec2c788,
32'h3e7300fa,
32'hbef57eb8,
32'hbb9a5d4a,
32'hbe455c37,
32'hbd3b1214,
32'h3f1260a9,
32'hbdba92c1,
32'h3cc01ae1,
32'hbf63ef9a,
32'h3ecfbdb6,
32'hbee12df2,
32'hbe353247,
32'hbe951a25,
32'h3e22bf5f,
32'hbe8a8516,
32'hbe88b2a7,
32'hbc5e0074,
32'hbb0431a5,
32'h3e2627f6,
32'hbea4060e,
32'hbd924e82,
32'hbefc12b2,
32'hbfb61147,
32'h3d1f6e49,
32'hbdcce050,
32'hbe8bc6ef,
32'h3eb64c59,
32'hbd5f3d33,
32'hbd59f4a5,
32'h3e65649e,
32'h3ea291b4,
32'hbed4c54f,
32'h3e42fe7b,
32'h3e228bf7,
32'hbcaecaae,
32'h3d8d4310,
32'hbdd6c4cc,
32'hbf138e4f,
32'hbf7d59e3,
32'h3ef9ae80,
32'hbe90a469,
32'h3e82a2e0,
32'hbd008709,
32'h3f413bf6,
32'hbf3c52ed,
32'h3d5a240c,
32'h3e1896a4,
32'hbce3ca56,
32'h3ec0546b,
32'hbf1d604f,
32'hbbe4c279,
32'hbf67a6f7,
32'hbe826a29,
32'h3dad29a5,
32'h3cfb6e33,
32'hbec2fff9,
32'h3e9b9c42,
32'h3ee1bba3,
32'hbdb23ba5,
32'h3c4eb73d,
32'hbc62e441,
32'hbf567b2f,
32'h3ed3760e,
32'h3d96eac5,
32'hbdbdbc2e,
32'hbe562ef4,
32'hbdf02d9e,
32'hbe985c2c,
32'h3e33fee2,
32'h3f08f5e0,
32'hbc763bd3,
32'h3e1cc3bb,
32'h3c085bf2,
32'h3e801d74,
32'hbdb1b6a5,
32'h3f12f432,
32'h3da33895,
32'hbe59731d,
32'h3f20e664,
32'hbf251bde,
32'hbe7cbc0b,
32'hbfc16896,
32'hbec60bc8,
32'h3d80363e,
32'h3d87f828,
32'hbedf3a9e,
32'h3d121820,
32'h3e2a47ed,
32'hbe65c7ca,
32'hbd7fd136,
32'hbe034e96,
32'hbe65b655,
32'h3f332826,
32'h3ec82bd4,
32'hbe9d1265,
32'hbe9192b5,
32'hbeab9d1c,
32'hbe628e37,
32'hbeda13ed,
32'h3eb302d3,
32'h3de7beb8,
32'hbf23a57a,
32'h3ef33787,
32'h3e0296fa,
32'h3e70f9c9,
32'hbed14d7e,
32'hbeb43cfb,
32'h3e1e9e40,
32'h3ee82f69,
32'hbf253d77,
32'hbf044ef4,
32'hbf24d631,
32'h3e0c5192,
32'hbd8049bf,
32'hbb48f01d,
32'h3b671553,
32'hbf75d9d7,
32'hbed19678,
32'hbe80261b,
32'h3d535fc8,
32'hbe82b06e,
32'hbe075673,
32'h3e11b66b,
32'h3ea14e9e,
32'hbe6896ad,
32'hbebb262c,
32'hbe782a41,
32'hbf96af8e,
32'hbe456ae6,
32'h3d0f170e,
32'hbdbc9990,
32'hbf3b6b4c,
32'h3ed5c792,
32'hbee5b615,
32'h3f5121c3,
32'hbde10aa4,
32'hbfcc604b,
32'hbe448c35,
32'h3da676ee,
32'h3e236e9e,
32'hbee6090c,
32'h3f1f86de,
32'hbd777c76,
32'hbd8e41c5,
32'h3d52f8ab,
32'hbf35c17d,
32'h3f65747d,
32'hbf015d03,
32'hbd2db877,
32'hbec1283f,
32'hbdd0bdc2,
32'h3eb65829,
32'h3f7f29d3,
32'h3e71a560,
32'hbe1867ee,
32'hbf432014,
32'hbef626f1,
32'hbf72e970,
32'hbea59d01,
32'hbe462e85,
32'h3f2515d0,
32'h3edcf703,
32'hbf0c03da,
32'hbe47088b,
32'h3f16ca84,
32'hbf0679a3,
32'hbfbba139,
32'h3e90cdde,
32'h3f207f62,
32'h3d59e1bd,
32'h3f1a90a6,
32'hbd43e4fc,
32'hbd2dbf8d,
32'hbc1ed824,
32'hbd676de9,
32'h3e95944b,
32'hbde16601,
32'hbda9193e,
32'hbf58bb0f,
32'hbf1d1796,
32'hbed7249b,
32'h3f11d054,
32'h3eb7d102,
32'hbfbfa447,
32'h3ee69796,
32'hbf203f06,
32'h3c520061,
32'hbd924613,
32'hbe5b4e30,
32'h3f3a05bb,
32'h3f5eb187,
32'hbd9b5486,
32'hbf2bdc0f,
32'hbdc8ffbe,
32'h3ea53920,
32'hbe54eece,
32'hbf41ebd7,
32'hbb09e682,
32'h3e2ee5ea,
32'h3de0914c,
32'h3e8863c3,
32'h3c15f021,
32'h3cf21277,
32'hbca23aed,
32'h3c7d70b1,
32'h3f45b752,
32'hbe49166b,
32'hbda05156,
32'hbf2af90c,
32'hbf0633e0,
32'hbc18f6bf,
32'hbe50a167,
32'h3cad14b9,
32'h3e3a0977,
32'h3db3e35d,
32'h3e0ee509,
32'h3f30b609,
32'hbe364f78,
32'hbcd7794d,
32'hbecbff8f,
32'h3eacf810,
32'h3d5fe8ab,
32'h3ebd660e,
32'hbcbcccac,
32'hbdc72182,
32'hbd65cd0a,
32'hbdbd9c65,
32'h3d23d6c7,
32'h3c8458b3,
32'hbd92f500,
32'hbd962e09,
32'h3dc02fe6,
32'hbc947d24,
32'h3d862aa0,
32'hbcda2c6c,
32'hbc5d3243,
32'hbb4755e7,
32'h3dd7a1d1,
32'hbb2351fa,
32'hbb61689e,
32'hbc844ce2,
32'h3c884b72,
32'hbd9350dd,
32'h3d30798c,
32'hbb9c182c,
32'hbd1e79db,
32'h3d12f812,
32'h3cbf7643,
32'h3da6c3dd,
32'hbd5f1a4c,
32'hbd4fd362,
32'h3c36554a,
32'hbb6dd509,
32'h3c813749,
32'h3c0cf324,
32'h3d28eb7e,
32'h3de04434,
32'hbc94b116,
32'hbae534d7,
32'h3d92b9f3,
32'h3dd1a988,
32'h3d06de23,
32'h3d31d1ca,
32'h3d264c0b,
32'hbdc5d2eb,
32'h3d6c44c8,
32'h3c248c2a,
32'hbbc0929d,
32'h3ca977ab,
32'h3c79d844,
32'h3d9c6bdf,
32'h3cf89eff,
32'h3bf85dc0,
32'hbe348ca1,
32'h3e297cb2,
32'h3b4940e4,
32'hbf200111,
32'h3f15ef39,
32'hbd0251b0,
32'h3ef01835,
32'h3d0e84ef,
32'h3d47a0a6,
32'hbc8e5a72,
32'hbdbc53f6,
32'h3d9c5aa5,
32'h3bdd88d0,
32'hbef87e8f,
32'h3dcf08d2,
32'h3f104eb9,
32'h3f9b2aea,
32'h3e7ee29b,
32'h3c0382ff,
32'h3ec04bdc,
32'h3d1f31da,
32'h3c88bb31,
32'hbf0c4f5e,
32'h3e5653da,
32'h3f092f00,
32'hbebe9c7e,
32'h3e43ca5b,
32'hbe1d3834,
32'h3eb6803e,
32'h3ece8878,
32'h3bdbbb64,
32'hbda1e4fb,
32'hbda07163,
32'hbed42445,
32'h3f269679,
32'h3eb82cf3,
32'h3e092112,
32'h3e98ab5c,
32'h3efc1b32,
32'hbdd0bf10,
32'h3f0802e7,
32'h3f20b9f9,
32'hbf577d5d,
32'hbf7310a3,
32'h3ed46df6,
32'h3e6da7cd,
32'h3f1daeed,
32'h3ee051e4,
32'hbeb2af63,
32'hbe47fca7,
32'h3dba67a9,
32'h3d55bc4b,
32'hbe5520a3,
32'hbf1669ee,
32'hbf404f10,
32'h3e0872b3,
32'h3eaf027c,
32'h3e55f183,
32'h3fad3c8f,
32'h3f175d92,
32'hbe6f297e,
32'h3ed778b6,
32'hbe1c0a84,
32'hbdb168cc,
32'h3ddc3986,
32'h3fad5576,
32'h3ea37fdf,
32'h3eeb0150,
32'h3ec439d1,
32'hbeab9b73,
32'h3f0b45cc,
32'h3f192f89,
32'h3d1c6c0a,
32'h3ebd4847,
32'h3ebcfa24,
32'hbed48bb4,
32'h3ecbb969,
32'h3f656f7a,
32'h3ee3fad2,
32'hbd37a0e5,
32'h3cb17eaf,
32'h3cb82f86,
32'hbf3831e0,
32'h3f0239e4,
32'hbe62418a,
32'hbf56f44f,
32'h3f29f7d5,
32'hbefce43b,
32'hbefa7bce,
32'h3e2e0e02,
32'h3e1b27b0,
32'h3e96514b,
32'hbe1aab32,
32'h3d7b140e,
32'hbe8307db,
32'h3f21526a,
32'h3e3d6c22,
32'h3db6f4b0,
32'h3df5345e,
32'h3d52543e,
32'h3b962b09,
32'h3f14aa1b,
32'hbe656701,
32'h3e11ca6c,
32'hbd777092,
32'hbf96e938,
32'h3f0dd699,
32'hbe178e71,
32'hbde78f3c,
32'hbf2c7c6f,
32'h3db4b79b,
32'hbbd7bf65,
32'hbeb8c36a,
32'h3e106625,
32'hbe546cb5,
32'hbe8e0738,
32'hbec38481,
32'h3e94fd5e,
32'hbe44d601,
32'h3ec9af3c,
32'h3f459f46,
32'h3e69870b,
32'hbf808d09,
32'hbd44075a,
32'hbe84a015,
32'h3f78b564,
32'hbed423c6,
32'hbcc81a94,
32'hbdbe08b5,
32'h3ee084b8,
32'hbf15f621,
32'hbe11ef0e,
32'h3d82f59b,
32'hbdabf4d7,
32'h3e28d75f,
32'hbe422b80,
32'h3ead939b,
32'hbec24cfe,
32'h3e33fab0,
32'hbebbbc0d,
32'hbb30aa2a,
32'h3c98d184,
32'h3cbf5333,
32'h3df59a9b,
32'hbeb9ef3b,
32'hbd82adfd,
32'hbcf20b3b,
32'h3e0f6174,
32'h3e6ec1ba,
32'h3c5aaf09,
32'hbd5fb5ac,
32'h3e6fa467,
32'hbf931aab,
32'hbe8e1926,
32'hbdf385b7,
32'h3eabebc9,
32'hbef4aaf5,
32'hbeccefbe,
32'h3edf9f9a,
32'h3d3704f5,
32'h3d68b506,
32'h3c25c310,
32'h3d063d6a,
32'h3db80dd2,
32'h3ee61bbe,
32'hbf3703e3,
32'h3ead03d8,
32'hbcdd7dae,
32'h3e8418b2,
32'hbf58404c,
32'hbc84d43c,
32'h3c4dfa7f,
32'h3d0a260a,
32'hbe0dcd8f,
32'hbf0400f1,
32'hbe3263af,
32'h3ceefd2a,
32'h3c789722,
32'h3ebcf715,
32'hbd9bfacf,
32'h3c2fd47c,
32'hbd731542,
32'hbf00cd77,
32'h3e8b2748,
32'h3d0a776a,
32'h3e69897b,
32'hbd236769,
32'hbf1b0898,
32'h3e2da8f5,
32'h3d162e05,
32'hbec2bf89,
32'h3a0ff815,
32'h3e334b58,
32'hbe33d3aa,
32'h3ed34710,
32'hbeb911d1,
32'h3e508817,
32'h3e357601,
32'hbd5a53e5,
32'hbebc4c25,
32'h3db64267,
32'hbcfcf006,
32'h3de21ed0,
32'h3d28b6da,
32'hbdcda700,
32'hbd535276,
32'h3e8902dd,
32'h3d93d1de,
32'hbcd1d18f,
32'h3e69cc02,
32'hbe942f6a,
32'h3e850cf3,
32'h3da39fe5,
32'hbd7e8f09,
32'hbe2ed8ef,
32'h3e8029e7,
32'h3eab801f,
32'hbf3ec9f4,
32'hbea2992d,
32'hbeb56c97,
32'h3ed77139,
32'hbf502df1,
32'h3eae6e57,
32'hbf062ed2,
32'h3db307ba,
32'hbedbe523,
32'h3e86c261,
32'hbda5d27a,
32'h3d2aed05,
32'hbeed5b97,
32'hbdcafdce,
32'hbca304ea,
32'hbe5bbcec,
32'h3d43b930,
32'hbd2b0915,
32'hbdbe3463,
32'h3dfdc87a,
32'h3ebfec46,
32'h3dda310c,
32'h3e41429a,
32'h3e665834,
32'hbd412c9d,
32'h3ea27851,
32'hbe676811,
32'h3e846bbc,
32'h3edd5feb,
32'hbd79edbf,
32'hbec38827,
32'hbddadfd5,
32'hbe674a0b,
32'h3e8a9ce9,
32'hbf1d3916,
32'h3d794f02,
32'hbdab92ca,
32'h3dac14e1,
32'h3d251d87,
32'h3d174fc4,
32'h3ea15f51,
32'h3e003622,
32'hbf69745f,
32'hbc9a6c60,
32'h3d4ac16f,
32'hbdeac50f,
32'hbe0528fa,
32'hbe2d8055,
32'h3e53612f,
32'hbdffcd60,
32'hbe956f20,
32'hbe44b2b6,
32'hbd61282a,
32'hbedb4338,
32'h3eae44ad,
32'h3e14bbf7,
32'h3d310e00,
32'h3e0d450a,
32'hbdcf262f,
32'h3e66aba5,
32'hbe082c67,
32'hbe216448,
32'hbf2c6626,
32'h3e6f1798,
32'h3d0dc135,
32'h3d70bc7b,
32'h3c9c0ae5,
32'h3ecd55c7,
32'h3e851ac5,
32'h3e1574d0,
32'h3da2e969,
32'h3ef4d105,
32'hbe5669a5,
32'hbd2210ea,
32'hbd2d76bb,
32'h3ca2c501,
32'h3e34640e,
32'hbbdb1b7b,
32'h3e6843e2,
32'hbea6425b,
32'hbe433dc1,
32'h3da30ce0,
32'hbdd41724,
32'hbf2cc7f3,
32'h3cb0b7bf,
32'hbe36bde4,
32'hbdeee0e9,
32'h3cd7fc42,
32'h3e37f268,
32'hbc32674b,
32'hbe23ecf4,
32'hbe2f7023,
32'hbf24fec6,
32'hbf6dc8a2,
32'h3db79226,
32'h3df2ffd3,
32'h3c7d2500,
32'h3eb04065,
32'hbdd60695,
32'h3ddc25ee,
32'h3e85bad5,
32'h3e6dcf51,
32'hbc96554a,
32'hbca4c1c9,
32'hbd48e8f7,
32'hbcbb3105,
32'h3b04d120,
32'hbd96529c,
32'hbe0c969e,
32'hbd6a7d5a,
32'hbeb6a5ef,
32'hbb96d2dd,
32'hbeb3dfb6,
32'hbe65fd5b,
32'h3d04597f,
32'hbca78e83,
32'hbe310c5f,
32'hbe441d76,
32'h3ecdd18c,
32'h3cfe611b,
32'h3e36e66b,
32'h3e0ff012,
32'hbec5e26d,
32'hbf95e1a2,
32'hbe098234,
32'h3d1558d2,
32'h3db7316d,
32'h3d01f984,
32'hbe3d0058,
32'h3e71c147,
32'h3e4e9591,
32'h3e18050d,
32'hbe253b2e,
32'hbaabd18e,
32'hbd237f24,
32'h3d83800e,
32'h3e2923aa,
32'hbdd1210d,
32'hbe023698,
32'hbda6cb61,
32'hbed2a29c,
32'hbd04ec48,
32'hbe2fdfce,
32'hbe63e49f,
32'hbca1eadb,
32'hbf13d8e9,
32'h3c4924ec,
32'hbd8e283e,
32'hbe826eec,
32'hbbb87cfe,
32'h3e624421,
32'h3d00b3c5,
32'hbea4a2e2,
32'hbea2dd66,
32'hbe2331eb,
32'h3d292673,
32'h3e8622bd,
32'h3cf66ab7,
32'hbd9f58fb,
32'h3e4e5c8e,
32'h3c4c8946,
32'h3d08a5e5,
32'hbdd4a5f0,
32'hbd965b18,
32'hbd5f0f42,
32'hbe86b23d,
32'h3e0d00f1,
32'hbe379410,
32'hbdea4905,
32'hbe14d245,
32'hbf2e6c07,
32'h3dc87e4e,
32'h3e3535a4,
32'hbe09c640,
32'h3c854953,
32'hbd5a3019,
32'hbe81abd5,
32'hbd9784af,
32'hbf0e1cb3,
32'h3d6e3848,
32'h3da08876,
32'hbdfb8d38,
32'hbf12bb29,
32'hbed2de67,
32'hbe4b7dc3,
32'h3cb33247,
32'hbc419900,
32'hbe454605,
32'hbe95a335,
32'hbcf5f2cd,
32'h3c95f352,
32'hbe7c07a5,
32'h3d55f715,
32'hbc96cf7f,
32'h3bab4e0f,
32'hbe994189,
32'h3e424b77,
32'hbda78131,
32'hbd9bb15a,
32'hbe8a21af,
32'hbfde4dee,
32'hbd0d8bd7,
32'hbee8ca7d,
32'hbe596471,
32'hbdd0f812,
32'hbe5eeeeb,
32'hbd9b008c,
32'h3d455392,
32'hbe23209f,
32'h3e5e58df,
32'hbe929f7f,
32'h3e116b12,
32'hbef822ab,
32'hbe28b3f6,
32'hbeb4a0da,
32'h3e3da5da,
32'hbe367db3,
32'hbe488681,
32'hbe060cf8,
32'hbe934224,
32'h3e9b129d,
32'hbdbee854,
32'hbe866932,
32'hbd5d1e7e,
32'hbd9b5646,
32'hbeae5772,
32'h3e0c3568,
32'h3cae834b,
32'hbd9a9b11,
32'hbd8703a7,
32'hbe6f7184,
32'hbd76f92e,
32'hbec33293,
32'h3d21d7a1,
32'h3e11cab8,
32'hbf1db6c2,
32'h3d17e9e1,
32'h3e1092e9,
32'hbd014abd,
32'h3e5c3ee4,
32'hbea905ed,
32'h3e546002,
32'hbee9411a,
32'hbe1bd26e,
32'h3e7c30f6,
32'h3d6c4eb6,
32'hbd47e0de,
32'hba54a318,
32'h3e4c17fb,
32'hbd98bd42,
32'h3c9bba59,
32'h3ebd5904,
32'hbed683e4,
32'h3bb97f09,
32'hbda250e6,
32'hbf0e7dd1,
32'h3d3eaa84,
32'h3db424a2,
32'hbcb87a89,
32'h3df2483b,
32'h3d86c598,
32'h3f0f10ff,
32'hbeb0bd18,
32'hbe1922ea,
32'h3e402df5,
32'hbe286e03,
32'hbea9e616,
32'hbdc1a7ed,
32'hbd456cab,
32'h3e05b1f1,
32'hbdc698cf,
32'h3da82764,
32'hbee9d9e9,
32'hbe0329fc,
32'h3ecc28cc,
32'hbe084e16,
32'h3e08fbc9,
32'h3cfdbeec,
32'h3e7256d3,
32'h3d05f36e,
32'h3cadfe72,
32'h3e1670b4,
32'hbdd8301f,
32'hbdb02838,
32'hbd0dfbe2,
32'hbe9994fc,
32'h3e6a70a7,
32'h3db6ad18,
32'hbd220065,
32'h3edefc05,
32'h3dbcb526,
32'h3eacfa88,
32'hbef833f7,
32'hbeff9e72,
32'h3c1335c1,
32'h3de07423,
32'hbebd1630,
32'h3e5b8881,
32'hbe68ecf1,
32'h3e7de9b3,
32'hbd8cf76b,
32'h3ddd8fd5,
32'hbefba76c,
32'hbc6e601c,
32'h3d1e69e2,
32'hbe124b39,
32'hbe9f13fd,
32'h3e6d4be4,
32'h3e3e248c,
32'hbe12d9d0,
32'h3e325821,
32'h3ef259e2,
32'hbef14aa3,
32'h3b83cd78,
32'hbdf71f92,
32'hbe232c8e,
32'hbddc361f,
32'h3e62d3d6,
32'hbe96c6f3,
32'h3d91f12a,
32'h3e3470a9,
32'hbe0fa264,
32'hbedb99d5,
32'hbf1e1d30,
32'hbbd7d018,
32'h3e6d81e4,
32'hbd8227be,
32'hbcda57d6,
32'hbd9c7c0c,
32'h3e560cdb,
32'h3d0fb639,
32'h3cff2c48,
32'hbd828aa2,
32'hbe3a24ee,
32'hbe1cad30,
32'hbf059c43,
32'hbeb73b53,
32'h3e3635e8,
32'h3d93030e,
32'hbd9d9052,
32'h3e3a6e97,
32'h3dc29b73,
32'hbfc6c356,
32'hbcfeccc5,
32'hbc80a160,
32'hbde3e0ce,
32'hbe99cae8,
32'h3e240ab8,
32'hbd95e81d,
32'h3db12645,
32'h3de7a56b,
32'hbe9bf17b,
32'h3c1c46ba,
32'h3dc8e0e8,
32'h3e3773fb,
32'h3ebcd839,
32'hbe33d1b2,
32'hbe147463,
32'hbe53ebfe,
32'h3e870b1b,
32'h3d897317,
32'hbe5aecf3,
32'hbe988838,
32'hbe415987,
32'h3e15e90c,
32'h3d57f61f,
32'hbc28b131,
32'hbda65a9a,
32'h3e4a654c,
32'h3e649c8c,
32'hbce2b2ae,
32'hbeb3b48a,
32'h3dab6e1e,
32'hbddc1fdd,
32'hbc6e585c,
32'h3c1f3a1d,
32'hbe93f0a4,
32'h3e26ed1a,
32'hbc82f7d0,
32'hbd188295,
32'hbd51c45e,
32'h3e150918,
32'h3cf63d01,
32'hbe0123f0,
32'h3cda09c2,
32'hbf34d3bb,
32'hbe51cf36,
32'hbec1abfd,
32'h3dafa559,
32'h3e759e6f,
32'h3ea4c43e,
32'h3eb46402,
32'h3e0df1f3,
32'h3d5f1fc5,
32'h3eaa5e25,
32'h3ec04218,
32'h3ec47814,
32'hbe334784,
32'h3dc66567,
32'hbe9b280d,
32'hbd2dd5dc,
32'hbf80e910,
32'hbf325e38,
32'h3d614b02,
32'hbd08baeb,
32'hbe8f6958,
32'h3e7e701f,
32'hbdf282ba,
32'hbe5102c8,
32'hbe893335,
32'h3e816705,
32'hbec55b74,
32'h3cfa1869,
32'h3dc0888c,
32'hbd1cdeba,
32'h3e3fba9d,
32'hbe38c490,
32'hbe01d636,
32'hbf4d3251,
32'h3d6371ef,
32'h3ea0d48a,
32'h3ebb25b2,
32'h3e87d9ad,
32'hbe83f7ed,
32'hbe430c39,
32'h3c288248,
32'h3e44a9ad,
32'h3da08517,
32'h3efb2a5e,
32'hbfc781aa,
32'hbe14dee1,
32'hbffa142c,
32'hbef26e5e,
32'hbd982eb9,
32'h3dafe2bd,
32'hbf719159,
32'hbf07bf28,
32'hbee8d304,
32'hbdfdfde9,
32'hbe19f039,
32'h3e8b43b8,
32'hbf71f741,
32'h3ebb8e18,
32'h3ef4a2b4,
32'h3ca48cff,
32'hbd0295d1,
32'hbe0ec415,
32'hbea92a68,
32'hbf090326,
32'h3e248329,
32'h3da037ee,
32'hbf5b8969,
32'h3d7d12db,
32'hbefdaf76,
32'h3dca92ac,
32'hbe5da37d,
32'hbf0464a1,
32'h3d2af1bb,
32'h3eb1d6c1,
32'hc0287cd8,
32'h3ec760ec,
32'hbfcd3541,
32'hbebbffba,
32'hbdbbfcc1,
32'h3cafd6ab,
32'hbfac3ab6,
32'hc00da28a,
32'hbf78291c,
32'hbe4374b1,
32'h3e63aab1,
32'hbf33cf41,
32'hbf04b867,
32'h3ead1c6f,
32'h3ea0530f,
32'hba288084,
32'hbd6e4188,
32'hbea26d32,
32'hbf278e86,
32'hbcd24c15,
32'h3ebb3c1e,
32'h3e34ebe1,
32'hbf90d979,
32'hbf1b5922,
32'hbf14e102,
32'h3e911934,
32'hbff26f7c,
32'hbfe5d6bd,
32'hbf9d1769,
32'h3f61b720,
32'hbf8cc633,
32'hbd894f45,
32'hbeceaebd,
32'h3eb69f16,
32'h3d3e2fdd,
32'h3d84580d,
32'hbf63683a,
32'hbe949c16,
32'hc0192fb8,
32'hbe3a493d,
32'hbf394f3d,
32'hbe846870,
32'hbd988d36,
32'h3e878bd6,
32'hbeda9648,
32'h3e319fc1,
32'hbf4b9cf9,
32'h3e8e1fbd,
32'hbfa61925,
32'hbe9bf6d1,
32'h3f304974,
32'h3e00a785,
32'hbe984292,
32'hbf1a13a8,
32'hbf01091e,
32'hbf1d19fe,
32'hbdd480a8,
32'hbfc5fb61,
32'h3e53b4e0,
32'h3f776cf6,
32'hbe0fca89,
32'h3e1731f4,
32'h3c2eb0ca,
32'h3e5cb3b3,
32'hbac9125b,
32'h3d79075d,
32'h3f25d0c9,
32'h3e1b153e,
32'hbe870401,
32'h3e7d1fe9,
32'hbb0dcccc,
32'hbdccedb8,
32'hbec448e0,
32'hbc662804,
32'h3fd1567f,
32'hbeb6f8e6,
32'hbf210fe9,
32'hbf5d012c,
32'hbef2639e,
32'hbf0c575f,
32'h3ea1da38,
32'h3ee61e9c,
32'hbd40d635,
32'hc0034476,
32'hbf0ac150,
32'hbed139a7,
32'h3e90b2e2,
32'hbf412502,
32'hbf6af9b0,
32'h3ded9fea,
32'h3d4bae13,
32'hbea5b5cc,
32'hbca3fa88,
32'h3ec69ee5,
32'h3c863892,
32'h3b3ffbc0,
32'hbe44679c,
32'h3e3cfe76,
32'hbe36259e,
32'h3fa0b747,
32'hbbb6e527,
32'h3e895fa0,
32'hbf59ce83,
32'hbf967317,
32'h3f3e82ad,
32'h3fba00d4,
32'hbe563197,
32'h3ed8dc7f,
32'hbec0fda5,
32'h3daa817a,
32'h3e230c8e,
32'h3f73ebfa,
32'h3c352821,
32'hbf691703,
32'hbd8d9da6,
32'hbc8b1ae6,
32'hbc82925c,
32'h3cee90cc,
32'hbc07ee7e,
32'hbd0c700b,
32'hbd485f7d,
32'h3d9e6bf9,
32'h3dae8f50,
32'hbd09196e,
32'hbd1c62a3,
32'hbb94375a,
32'h3bbcd442,
32'h3d0eb773,
32'h3c1e015a,
32'h3c801aa1,
32'h3b5dd517,
32'hbd4190e5,
32'h3d7ad107,
32'h3d1769ac,
32'hbdac073d,
32'hbd9f85f6,
32'hbd22739d,
32'hbcbb0f37,
32'h3db02441,
32'hbdc12cd9,
32'hbd0850fc,
32'hbcfedca5,
32'h3d039436,
32'h3d64d041,
32'hbca9fa79,
32'h3ee64c19,
32'h3e7e5b02,
32'h3db9ef0c,
32'h3ea6c185,
32'hbd8837be,
32'h3fbf79eb,
32'h3fd7b4e8,
32'h3d50cc33,
32'hbd41dbfb,
32'h3cca502a,
32'hbd6e4bc6,
32'hbf17d8d7,
32'h3de4c4c1,
32'hbd4c6643,
32'hbfa65216,
32'hbd43f9df,
32'hbdc3c777,
32'h3dd092e2,
32'h3e5cb8cf,
32'hbeee0214,
32'h3e21e808,
32'hbd9ffb00,
32'hbfe85a3e,
32'h3fabdb79,
32'h3fd47f7f,
32'h3f0a77ef,
32'h3e84b274,
32'h3d126d01,
32'hbef682a6,
32'h3d888333,
32'h3f1ac2ec,
32'hbdb03015,
32'hbf09f8de,
32'h3eb4adf1,
32'h3ed17cec,
32'hbe675eba,
32'h3e8715cd,
32'hbdd0e31d,
32'h3f2d031f,
32'h3c38dac6,
32'h3de6278b,
32'h3fbe14e9,
32'h40080847,
32'h3fbab7b9,
32'hbf155307,
32'h3e0d6cfc,
32'hbe3a17fa,
32'h3ed45f69,
32'h3f3c723b,
32'h3db1e974,
32'hbd9e0d43,
32'h3d5be843,
32'hbf6b2d30,
32'hbe8e2977,
32'h3f628cf0,
32'hbe7092f6,
32'h3ed75c74,
32'h3f27f8f5,
32'hbed7528e,
32'h3f0d159f,
32'h3f736866,
32'h3f4ed0fa,
32'hbf17a91e,
32'h3f30393d,
32'hbb109346,
32'h3f370ec3,
32'h3f8613e7,
32'h3f22a450,
32'h3ebf8985,
32'h3ccf80ec,
32'hbac67825,
32'h3da922ac,
32'hbf7adc17,
32'hbebcc80a,
32'hbe79deae,
32'hbf465626,
32'h3dc04f3d,
32'h3fa744c4,
32'h3cfa2540,
32'h3e054d3d,
32'h3e38b72d,
32'hbb8427e7,
32'hbf883d59,
32'hbf0ed944,
32'h400770ff,
32'h3eebf8b1,
32'h3f198114,
32'h3eb76ec8,
32'hbe585e31,
32'h3f2472b5,
32'h3d8de354,
32'h3df79a74,
32'h3eecd958,
32'hbe8b17bb,
32'hbf67e915,
32'h3f0db25e,
32'h3f0ad43d,
32'h3f09e123,
32'hbe17ac64,
32'hbb4033f8,
32'h3d4f605d,
32'hbf8030f4,
32'h3ed041c6,
32'h3ec489cf,
32'h3e64086c,
32'hbeab9e3b,
32'hbed15dcb,
32'hbee35668,
32'hbd686842,
32'h3f0961a4,
32'h3e7a7a82,
32'hbe8e3516,
32'hbec73b29,
32'hbf041adf,
32'h3e3d3459,
32'h3f1ebe73,
32'h3d0ebbc8,
32'hbd36624c,
32'h3f4aeb85,
32'h3e096c6f,
32'hbe83c0a6,
32'hba455f55,
32'h3efce526,
32'hbeec1fbc,
32'hbf0a2644,
32'h3eb35439,
32'h3d92dc9f,
32'h3d8690bb,
32'hbf7ddb1c,
32'hbd904b28,
32'hbd727a58,
32'hbf1fa722,
32'hbe15ba53,
32'h3f15f89e,
32'hbe39c689,
32'hbea92eca,
32'h3e896dc5,
32'hbe2581de,
32'h3e99d715,
32'h3ed63503,
32'h3eabd2ce,
32'hbf00ca3e,
32'hbd74bff7,
32'hbe1da1cf,
32'h3d30e05f,
32'hbe4bbb64,
32'hbf243fe3,
32'h3eb3f4c6,
32'h3e9582a3,
32'h3d3261ca,
32'h3e931c97,
32'h3de81ea2,
32'h3e98a03e,
32'hbdb152cb,
32'hbc84ea5b,
32'hbd8dcd37,
32'hbecbd6a7,
32'h3e6475d9,
32'hbec33c8f,
32'hbd315ba4,
32'hbc9283f5,
32'hbe36a3cd,
32'h3e94f336,
32'hbebeccd9,
32'hbd5a4cfd,
32'hbe8ce05b,
32'h3eb10627,
32'h3f15de38,
32'h3d8539cf,
32'hbe852e58,
32'h3ac873b5,
32'hbf8c9d13,
32'hbead0d1c,
32'h3d1ded17,
32'h3f0811d9,
32'hbe99948b,
32'hbe073352,
32'h3f456807,
32'hbd030dfd,
32'h3e12363b,
32'h3f68f5d8,
32'h3db34b06,
32'h3e176a6b,
32'h3ccc41f4,
32'hbeff49ed,
32'h3e151868,
32'hbea973d8,
32'h3e650756,
32'h3e592256,
32'h3d895eba,
32'h3d2ca199,
32'hbb46fbf7,
32'h3e7d8ce4,
32'hbe60d8c1,
32'hbdc83cc0,
32'h3d1f44c4,
32'h3d375496,
32'h3bdfaeaa,
32'h3d5047cd,
32'hbf03de0a,
32'hbc89be63,
32'hbe55348c,
32'hbc8108d7,
32'hbd6fa6ea,
32'h3ec094fa,
32'hbe3cfb37,
32'h3f1c7619,
32'h3f0a768f,
32'hbd80d3ea,
32'h3dd6740a,
32'h3e64a425,
32'hbe5f4346,
32'hbf02aa6b,
32'hbe902415,
32'hbeaa1fb4,
32'h3c81f635,
32'hbeddb86f,
32'h3e04ddfc,
32'hbe1527c7,
32'hbd242cc8,
32'h3c416dae,
32'hbe27eb5c,
32'h3e3d4ca0,
32'h3d09026a,
32'hbe0802d9,
32'h3e6d62a6,
32'h3de713ea,
32'hbeccf09b,
32'h3e277698,
32'h3e3a5959,
32'h3d98a876,
32'hbeff656f,
32'hbe25eb38,
32'h3dfd0d4f,
32'hbdbc7307,
32'h3ec9b88e,
32'h3d77892d,
32'h3eaa1d3b,
32'hbe91e1ec,
32'h3ecdc941,
32'hbd3732f6,
32'h3d8b1dfc,
32'hbe014224,
32'hbea300ee,
32'h3ddbfe47,
32'h3d7bcce6,
32'hbeb048c9,
32'hbc4a1f3f,
32'h3e4d3b64,
32'hbb133f36,
32'hbd418591,
32'hbe881b5a,
32'h3e296f16,
32'h3e21d495,
32'hbe5f22b8,
32'hbd5ab74b,
32'hbe80d634,
32'hbded90d4,
32'h3cc25904,
32'h3ebfb216,
32'hbe02fb9c,
32'hbd8f26f6,
32'hbe80a177,
32'h3ee8681a,
32'h3f431853,
32'h3e08ad7d,
32'hbe595852,
32'h3e09eade,
32'hbf5ad949,
32'hbe76be98,
32'hbeaea994,
32'h3d04cb6b,
32'h3ea24381,
32'h3d20d8bc,
32'h3efebef5,
32'hbddcc841,
32'hbd9f0a1c,
32'hbe915b82,
32'hbe364bf0,
32'hbd869a2c,
32'hbd8e2e41,
32'h3c18973c,
32'h3dddf45b,
32'h3cc85891,
32'hbc124d26,
32'h3b169ed8,
32'h3adafb30,
32'h3dd9ef78,
32'hbe724e57,
32'hbe88118e,
32'hbde073d4,
32'hbf423b89,
32'hbe22cb96,
32'hbd6e1edf,
32'h3f06406b,
32'hbe65927d,
32'hbd972624,
32'h3cbeb9d7,
32'hbf34ad71,
32'hbe773fa9,
32'hbec50aed,
32'hbdf6f9df,
32'h3e8297d1,
32'h3ea97ced,
32'h3e5cccae,
32'hbd9d3bf1,
32'hbf075a4a,
32'hbd4d8f8b,
32'h3c8452a4,
32'hbba69bac,
32'hbdadfd1a,
32'h3e624f19,
32'h3ec160f3,
32'h3dab2736,
32'h3d775ae3,
32'h3c70e39a,
32'h3e147974,
32'h3d8a9584,
32'hbe2e38e3,
32'hbe9068f8,
32'hbdeb668b,
32'hbeecc097,
32'h3df4a0fe,
32'h3eb25dc2,
32'h3e226d7a,
32'hbe027ef6,
32'hbe3877d0,
32'h3d710f31,
32'hbf07c77a,
32'hbeaf2844,
32'hbf1187b9,
32'hbded215d,
32'hbd92e6cf,
32'h3e3657cf,
32'h3ddba4cd,
32'h3e15511d,
32'hbe5dfc06,
32'hbda0b2ac,
32'h3eda505e,
32'h3d94d3f1,
32'hbadf8f4a,
32'hbe7735f7,
32'hbdaf4364,
32'h3d867d53,
32'h3dbb1293,
32'h3e37786d,
32'hbd7729c6,
32'h3e50c8a1,
32'hbecc7f9e,
32'hbf04c9c3,
32'h3bd15f64,
32'hbf1293d3,
32'hbda49a16,
32'h3e15bf92,
32'hbe1e2c45,
32'h3d363f2a,
32'h3e56b2b1,
32'hbe70f07c,
32'hbece1cee,
32'hbe8e0ff8,
32'hbedccb0e,
32'hbd5a224f,
32'h3c4bc56c,
32'h3e34279f,
32'hbe904047,
32'h3e8a43a3,
32'hbe37e44f,
32'h3e3ac4d9,
32'hbe72fa4d,
32'hbd9ff35f,
32'hbda21708,
32'hbe26b068,
32'h3e91e337,
32'h3c399780,
32'hbb15f3db,
32'h3e107813,
32'hbd253d30,
32'h3e18fa63,
32'h3c982924,
32'h3c8e6ba7,
32'h3e589535,
32'hbee59a58,
32'hbe05bd82,
32'h3e8eca1d,
32'hbe765338,
32'hbd8a525a,
32'hbcad193a,
32'hbe2dd66d,
32'hbbd03fc7,
32'h3c96b739,
32'hbe6e96ca,
32'h3d9e9071,
32'hbd8df5b0,
32'hbe5362c1,
32'hbd6cea5f,
32'h3e2f6008,
32'hbda23cf1,
32'hbd3be16b,
32'h3dc8b9e1,
32'h3caa094d,
32'h3da9aaaf,
32'hbe176ccf,
32'h3e2e96b1,
32'hbe579c44,
32'hbe9c8d3a,
32'hbd25c6d0,
32'hbf8e1a35,
32'h3e1e74cf,
32'hbe2aeadc,
32'hbe1df718,
32'h3d6c51a6,
32'hbddd30b4,
32'hbd19dfe8,
32'h3e713baf,
32'hbef55da3,
32'h3c66981a,
32'hbea13996,
32'hbd1ad535,
32'hbe9bcf13,
32'hbe8174bb,
32'hbe316b54,
32'h3d2c538c,
32'h3dc01c05,
32'hbe9d15fd,
32'hbea02463,
32'hbedca664,
32'h3ded5a9a,
32'hbe742ed1,
32'h3d2d9e42,
32'h3d3c01d4,
32'hbbbc1894,
32'hbe592a70,
32'h3e1122f0,
32'h3db5885a,
32'hbd0ffe51,
32'hbee006c1,
32'hbf90f601,
32'h3c216f6f,
32'hbeb1c4d5,
32'hbc8ba0ac,
32'h3ca1d27f,
32'hbdf0a55f,
32'hbd1a0b19,
32'hbe011b60,
32'hbf0f1e88,
32'h3d6f08f8,
32'hbefd2d9c,
32'h3d780029,
32'hbf07eef5,
32'h3d909c00,
32'hbe33406e,
32'h3dde7d79,
32'hbd02a61e,
32'hbe86516f,
32'h3d615c2b,
32'h3d87ef92,
32'hbbc18db9,
32'hbee56232,
32'hbd33fc4a,
32'hbe09cad8,
32'hbd8eda3f,
32'hbf263d7d,
32'h3e2fbeec,
32'hbe0ccdcc,
32'hbe1dfb9d,
32'hbdb8d340,
32'hbeea5bcc,
32'h3e8f260d,
32'hbe9d6d69,
32'hbe095e8a,
32'hbdd95fd6,
32'hbf16e131,
32'hbe48e64b,
32'hbe00b273,
32'hbe838ef8,
32'hbd1e0429,
32'hbe436729,
32'h3e7ad366,
32'hbe2391bf,
32'h3e1378e0,
32'hbe988cb0,
32'hbbeb917b,
32'h3ebf27ee,
32'hbedab920,
32'h3cdb2845,
32'h3dbba3e1,
32'hbe283e5f,
32'hbe1a60c3,
32'hbe7b5192,
32'hbbf660f3,
32'h3d2829aa,
32'hbed018bd,
32'h3d60cd11,
32'hbe693315,
32'hbe82c0e4,
32'h3e6fd16c,
32'hbd5b337e,
32'h3e8b8b7a,
32'hbe4fdba4,
32'hbe08786a,
32'hbd09eb24,
32'h3e60ff0e,
32'hbea4fd19,
32'h3e05b9b1,
32'h3d800bdf,
32'hbd0cccaa,
32'hbe8ec626,
32'h3db61eb7,
32'hbe1cedd7,
32'hbd71504f,
32'hbe5547aa,
32'hbd33f02e,
32'h3f137831,
32'h3cdf2716,
32'h3ed17112,
32'hbe86cc47,
32'hbe368fbc,
32'hbe8b578e,
32'hbd0ebd71,
32'hbdb1294d,
32'hbd1c2180,
32'hbe0620c4,
32'hbde0c2d7,
32'h3df8bc5e,
32'hbe14052c,
32'h3e307bec,
32'h3e5b4762,
32'hbdf3251c,
32'hbec4f85a,
32'hbed1118f,
32'hbcfff5e0,
32'hbdf62f1b,
32'hbe117eae,
32'h3d84b3b9,
32'hbda8bfe3,
32'h3dfb16ad,
32'hbdafc30d,
32'hbe82aeac,
32'hbefde395,
32'h3e209b52,
32'h3d78af05,
32'h3e385c34,
32'h3eb14d8c,
32'h3ddd1ba0,
32'h3d6fc31c,
32'hbcdb2ae6,
32'hbdaed417,
32'hbc073523,
32'hbe1efc60,
32'hbd8d06c2,
32'h3d135689,
32'hbde07496,
32'hbe92dfbb,
32'h3ebec126,
32'h3baabf1d,
32'h3e3a0420,
32'h3ea0876e,
32'h3d66a451,
32'hbd77f057,
32'hbe93e43e,
32'hbd59d57c,
32'hbee4a8f1,
32'hbe14d3b7,
32'hbce8fca9,
32'h3d1757f5,
32'hbda69459,
32'hbdb4363a,
32'hbc134049,
32'hbe91dda9,
32'hbe65b583,
32'hbe461638,
32'hbe80baaf,
32'hbe1dfb6b,
32'h3e1798e5,
32'h3deeaf5a,
32'hbe85dbd0,
32'hbd4d1138,
32'h3cd9c308,
32'hbf68e808,
32'h3b807af7,
32'h3d8985ec,
32'hbd2d9f80,
32'hbeadc6f0,
32'h3dd5d260,
32'h3e3a148e,
32'h3b884916,
32'h3ce0c06e,
32'h3e5e13f4,
32'h3e984e64,
32'h3e27923e,
32'hbdb5de0a,
32'hbf1d07dd,
32'hbe9b8776,
32'h3d99deb5,
32'hbea81f3f,
32'hbe1b878b,
32'h3e9c3fec,
32'h3daddb55,
32'hbc9b0640,
32'h3e4e2752,
32'hbeb764c6,
32'hbea4e139,
32'hbeef7220,
32'hbcb2ecee,
32'h3e3b0e9b,
32'hbe3dd3d5,
32'hbe60461e,
32'hbe583671,
32'hbec8908a,
32'hbd956145,
32'h3d89000c,
32'hbe5963d3,
32'hbe7db9fe,
32'h3ecda58a,
32'h3e225455,
32'h3dce7c2f,
32'hbe0083e9,
32'hbe070fce,
32'h3da259aa,
32'h3d538a2d,
32'h3e5f64b3,
32'hbeb0ebd8,
32'hbeab6ad3,
32'hbe960d4a,
32'hbe37b9a4,
32'hbc4266fd,
32'h3eb116e4,
32'h3d87b492,
32'h3e8dd22f,
32'hbe42c3f1,
32'hbf006870,
32'h3e0989e9,
32'hbd974b03,
32'hbdf10eb4,
32'h3e985c46,
32'hbea15a58,
32'h3e39db19,
32'h3e9f39c2,
32'hbee86774,
32'h3c963140,
32'hbd59afb3,
32'hbe510ca8,
32'h3ec35aee,
32'h3ebd074c,
32'hbca24887,
32'h3e278a5c,
32'h3ec7aafe,
32'hbccb9e6b,
32'h3ed02435,
32'h3d8af17b,
32'h3da8ced1,
32'hbf4a3d18,
32'hbec1287b,
32'h3d82f4b2,
32'h3d616257,
32'h3e819baf,
32'h3ef65cb4,
32'h3efdaa01,
32'h3eaa12ee,
32'hbe00f18a,
32'hbc9ce299,
32'hbf22d623,
32'h3da9fb61,
32'h3f0206fa,
32'h3ea352a1,
32'hbf761cd9,
32'h3e14f642,
32'hbf2056f6,
32'hbf87b1b5,
32'h3d41f0ad,
32'hbc6735f0,
32'hbf1c6646,
32'hbd929908,
32'hbe02f247,
32'h3e1a671a,
32'hbeeaeade,
32'h3ea28d4d,
32'hbf0d4576,
32'h3ea3b6d8,
32'h3ef79cac,
32'hbe832e41,
32'hbf1998c1,
32'hbeb6b74d,
32'hbee90da6,
32'h3ea6756e,
32'h3e55b109,
32'h3edd39b8,
32'hbf4405a9,
32'h3d5db680,
32'hbfd00daa,
32'hbea1d7d7,
32'hbf1ff081,
32'hbf281c10,
32'h3df89f7d,
32'h3f0496f0,
32'hc00c4309,
32'h3df38ab4,
32'hbfb9183a,
32'hbf5b32bd,
32'hbd96fb65,
32'h38f3fd5a,
32'hbf3831f0,
32'hbe5afede,
32'hbf050b70,
32'hbee2c020,
32'hbf31ec51,
32'hbeca7d2e,
32'hbf580fdc,
32'hbe5c5913,
32'h3ea460aa,
32'hbc2b02b0,
32'hbf99bb82,
32'hbe58f26d,
32'hbeb54735,
32'h3eb426de,
32'h3f2c4972,
32'h3e2a811f,
32'hbf624444,
32'hbf4657e3,
32'hc006b8e1,
32'hbf0e280d,
32'hbf85f4ee,
32'hbff391f2,
32'hbdd9a7e3,
32'h3f072315,
32'hbfaea710,
32'hbe91b1df,
32'hbeeb1f7e,
32'hbeb64ba2,
32'h3cda2ae6,
32'hbd045596,
32'hbef3beb8,
32'hbecb245f,
32'hbfb092fb,
32'hbedb8aa5,
32'hbf8c03a0,
32'hbeb468a4,
32'hbf0f84f8,
32'hbe82fe11,
32'hbe5820f9,
32'h3e22a2a9,
32'hbebb105a,
32'hbda28244,
32'hbf98484b,
32'hbf8fe876,
32'h3f4c7545,
32'h3d0f195d,
32'hbef5e265,
32'hbfb2c58e,
32'hbf4e7180,
32'hbf13c9bd,
32'h3e2e6af9,
32'hbfe14969,
32'h3eba76fe,
32'h3e5779bd,
32'hbe91fd35,
32'h3eb94f21,
32'h3c1b4f88,
32'h3e481acc,
32'hbcf51d52,
32'h3d20c0fb,
32'h3eeb3641,
32'h3e10360c,
32'hbeaa3bcc,
32'h3e4e45e7,
32'h3dbb60a3,
32'hbe5e406a,
32'hbeeb9642,
32'h3e93eb34,
32'h3f3b2982,
32'hbe3a425e,
32'hbf099381,
32'hbf00ed03,
32'hbedf738f,
32'hbea6e4ca,
32'hbd7335a4,
32'h3f31de4f,
32'h3bd8eac3,
32'hbfa62569,
32'h3e623e61,
32'hbf28a202,
32'h3dd825f2,
32'hbf2e3918,
32'hbf16cf2d,
32'h3f357d99,
32'h3df48aeb,
32'h3ea71d83,
32'hbda8cada,
32'h3e924c98,
32'h3d9b8329,
32'hbd3a09a7,
32'hbeb0ea07,
32'hbd998e30,
32'hbdc2142d,
32'h3ef6269c,
32'h3d4c4d9f,
32'h3e1d50f1,
32'hbe5867dd,
32'hbe9c0a06,
32'hbf391e55,
32'h3f63ca48,
32'hbc494ae1,
32'hbfc56bc6,
32'hbe2ac57a,
32'hbd3e2f86,
32'h3edf2ec0,
32'h3fba8e7e,
32'h3dca7234,
32'hbf4760d8,
32'h3da68499,
32'h3f0c89bf,
32'h3ea2beea,
32'h3e5eae51,
32'hbcc7de75,
32'h3d9de49d,
32'hbc073e81,
32'h3e1cde1b,
32'hbbcb1284,
32'h3d4686a8,
32'h3cb34ce0,
32'hbd44e280,
32'h3ee74353,
32'hbd85a8d2,
32'hbcdaa9b0,
32'hbee3b33a,
32'h3d48dd03,
32'h3d646515,
32'h3d0d791c,
32'h3e0b3bd7,
32'hbd934b50,
32'h3dc8af5e,
32'hbddc2346,
32'h3da9f0f4,
32'hbe0c24a9,
32'h3db6f2e7,
32'hbe856d85,
32'h3c6f8046,
32'hbc11660c,
32'h3e421875,
32'hbdde26ad,
32'h3fb868cf,
32'h3f8f92f8,
32'h3d1a4f07,
32'h3f5e9c81,
32'h3df21aa1,
32'h3f271e1d,
32'h3f9f3684,
32'h3fbaab86,
32'hbc83ee40,
32'h3d3198d4,
32'hbc01302e,
32'hbf3323ca,
32'h3eab5145,
32'h3f369122,
32'hbde8ac38,
32'h3c963e85,
32'hbe84c4e5,
32'h3f666082,
32'h3e8fdfc1,
32'hbf97ce48,
32'h3ea6f159,
32'hbde40577,
32'hc004d802,
32'hbee66266,
32'h4012ecee,
32'hbda9aa5c,
32'h3f4e3320,
32'hbd44d0f7,
32'hbfdf9094,
32'h3dce84d1,
32'h3f1ad7fe,
32'hbcfd89af,
32'h3e76e27a,
32'h3e864a60,
32'h3dd8b1cc,
32'hbf63e63e,
32'hbf3ccec5,
32'hbe81ca8a,
32'h3ef55570,
32'h3d2e5636,
32'h3dc23ef1,
32'h3e906bfd,
32'hbf96a42e,
32'h3e9f2eec,
32'hbf324fcf,
32'hbdbd5740,
32'h3e8b95e2,
32'h3f7fb946,
32'h3f097c3d,
32'h3ea0945c,
32'h3c3892dc,
32'hbbaa4dc6,
32'hbec8441c,
32'hbdeabe08,
32'h3fd18c4f,
32'hbef3dc65,
32'hbcc8d1d6,
32'hbe26274c,
32'h3e0cdde1,
32'h3f8602ae,
32'h3f10d43e,
32'h3f023d68,
32'hbdd4c3ed,
32'h3f4d5262,
32'hbdb0d27b,
32'h3d34f13a,
32'h3eadd10b,
32'hbf6f368e,
32'h3ebfc6ba,
32'h3d06719b,
32'h3d21ea55,
32'h3ed9facf,
32'hbf928ae8,
32'hbde19b6a,
32'hbe4d69ae,
32'hbf303798,
32'h3f06fa4f,
32'h3e96ef39,
32'h3e299d60,
32'hbd6aae75,
32'h3e9b05cd,
32'hbf357bb9,
32'hbed58ae6,
32'h3e0c5fec,
32'h3f632423,
32'h3e65816a,
32'hbd2069ab,
32'hbe42cd8f,
32'hbf1c1115,
32'h3f2db75a,
32'hbca7928d,
32'h3f07afcc,
32'hbd675477,
32'hbf158aed,
32'hbf2f2342,
32'h3f68ad06,
32'hbe17ba97,
32'hbeee29fb,
32'hbe1bca7d,
32'hbda1fa8e,
32'hbc6c8a29,
32'hbee921e9,
32'hbe3fb33b,
32'h3e8baa24,
32'h3e102505,
32'hbd155159,
32'h3f0114b1,
32'hbe918470,
32'h3c6d5510,
32'hbe146550,
32'hbe13e49b,
32'hbf69c869,
32'hbdb74904,
32'h3dfadf3f,
32'h3d3ccf24,
32'h3bb813b0,
32'h3cc700f0,
32'hbec6cd85,
32'hbf075d1d,
32'hbdd69bae,
32'hbc392bad,
32'hbe4a0612,
32'h3d1f862e,
32'hbf8a8876,
32'hbea148e1,
32'h3e4fa08d,
32'hbeb642ca,
32'hbf01fe0a,
32'hbba3449f,
32'h3bcd31c8,
32'hbcaf9ecb,
32'hbe5bd42b,
32'hbda3d5ca,
32'hbdd45ee0,
32'h3e2f413e,
32'h3dab3bc2,
32'h3ea9bbb4,
32'hbd72cd48,
32'h3d25aa67,
32'hbda53181,
32'h3da3a28f,
32'hbf95ce98,
32'hbbeb6d56,
32'hbeb83eda,
32'hbdc2cd88,
32'hbe54c26d,
32'hbf46f42f,
32'h3eb617eb,
32'h3f0a260c,
32'hbee95fad,
32'hbe86a129,
32'h3c6bc427,
32'h3e213fbc,
32'hbe844b0e,
32'hbeeb6c50,
32'h3e1b1269,
32'hbda72791,
32'hbe4a8463,
32'h3cfe6e12,
32'h3d4571d4,
32'h3d403bb7,
32'hbe25f089,
32'hbe6bce2f,
32'hbe772422,
32'h3e39fba1,
32'hbf11a2f9,
32'hbcbe7644,
32'h3e43776e,
32'hbdc8edb2,
32'hbdf6c982,
32'h3d95bfc2,
32'hbfd5f7bb,
32'hbee4308c,
32'hbe94cce4,
32'hbe04f769,
32'hbdce2cb5,
32'hbe06fede,
32'h3f18aa23,
32'h3edc702f,
32'h3e4527d0,
32'hbe6b89b4,
32'h3e817130,
32'hbcf00605,
32'h3c8c4e64,
32'hbe6eab30,
32'hbdb511f1,
32'hbf1af541,
32'h3e180cf8,
32'h3d8ec4b6,
32'hbcf89e8c,
32'hbc53334f,
32'h3db47c2b,
32'h3d92fe9c,
32'hbbcddef0,
32'h3dae793a,
32'hbe10e9b5,
32'h3d828010,
32'h3e7c549f,
32'hbdb13985,
32'h3e6e9a00,
32'hbd93325a,
32'hbe8cde34,
32'hbe84f56f,
32'h3d7c2024,
32'h3e5867f9,
32'h3e4e091d,
32'h3e0976d7,
32'h3e143ddd,
32'hbc63fd72,
32'h3d917df7,
32'h3df721cb,
32'h3dba830d,
32'h3d63c9aa,
32'h3e875daf,
32'hbe90c9db,
32'hbe80c664,
32'hbe1c19ee,
32'hbe00a474,
32'hbf62a346,
32'h3c992d2c,
32'h3c7fd7f8,
32'hbe49879d,
32'hbde7bc67,
32'h3e4ceec1,
32'h3db8b58c,
32'hbd8de0a8,
32'h3d8f852c,
32'h3e83cd6e,
32'hbdd78f52,
32'h3d4d06a4,
32'h3e12101d,
32'hbc93032b,
32'hbea97f6e,
32'h3d67098c,
32'h3cfde655,
32'h3bf6c0e1,
32'hbe0233bb,
32'h3d5c8bcb,
32'hbf14b24a,
32'h3d057814,
32'hbda73f70,
32'hbda9df48,
32'hbe1b1907,
32'h3d81edbf,
32'hbe0fa75f,
32'h3d5b335f,
32'hbf46fad3,
32'hbe2c695d,
32'hbf088a67,
32'hbd379e9f,
32'hbd9f0a0d,
32'hbd97aa5b,
32'h3e28ad49,
32'h3e20b469,
32'hbd073e6f,
32'h3eb33192,
32'h3df36c22,
32'h3cbac27f,
32'h3d2621c9,
32'h3e07fac0,
32'h3dfb636e,
32'hbe0382bf,
32'hbdf23b28,
32'h3e610eed,
32'h3e4c5f30,
32'hbe593291,
32'hbee2333d,
32'h3c351ce7,
32'hbef2fb60,
32'hbe406c21,
32'h3e233a26,
32'h3db0a03d,
32'hbeac3127,
32'hbe029324,
32'h3d98b0b9,
32'h3eb75aa6,
32'hbf58620d,
32'h3df64f54,
32'hbe3ab596,
32'hbe2285b1,
32'h3d88e9e0,
32'hbd92998b,
32'h3eec66f9,
32'hbd4ca613,
32'hbd542c53,
32'h3e5b33c3,
32'h3e05641d,
32'h3de816a5,
32'hbe2a0188,
32'hbe5cc76b,
32'hbe4d7860,
32'hbf3804b6,
32'hbdd3fc06,
32'h3e835bfc,
32'h3eddf5d4,
32'hbe22e3bb,
32'hbed1fd3d,
32'h3e383ce7,
32'hbecbc7ff,
32'hbf181f69,
32'hbd1bf010,
32'h3da71975,
32'hbdb57036,
32'h3d35e6c3,
32'h3ebef2df,
32'hbeb56bbc,
32'hbf8f724b,
32'h3ddd118b,
32'hbeab298c,
32'hbd02d70c,
32'hbcd8468c,
32'hbe942e57,
32'hbe008b5e,
32'hbd27be67,
32'h3d838905,
32'h3ed9be27,
32'h3c11fa22,
32'h3e8160b9,
32'hbdfdf89a,
32'hbe43de74,
32'hbdd13942,
32'hbee86c05,
32'h3d9b9903,
32'h3ee2662d,
32'hbbc06cfe,
32'hbdc1085e,
32'hbe5c278f,
32'h3db2ce83,
32'hbe95a25a,
32'hbf60657a,
32'h3da444c8,
32'h3d394914,
32'hbd664fb3,
32'h3c4077b2,
32'h3e7e5c56,
32'hbddca914,
32'hbec91b89,
32'hbdd32691,
32'hbe9c8110,
32'h3bc3bdf6,
32'hbd2f3924,
32'hbe5d64b7,
32'hbe6c4759,
32'hbe66cc0d,
32'hbc6720be,
32'hbd6baaa9,
32'h3e722306,
32'h3e475c24,
32'h3e3d0117,
32'hbdcce18f,
32'h3dbfd421,
32'hbe203bd1,
32'hbda6e4b1,
32'h3dd81fae,
32'h3d89fed7,
32'hb9fe9b41,
32'h3b238c76,
32'h3d9d86e2,
32'hbe501238,
32'hbf548f8d,
32'hbe5aeeea,
32'hbdf4af8f,
32'hbe135908,
32'h3e70b151,
32'h3d267bc3,
32'h3dd2ca57,
32'hbf2a0d1b,
32'h3e265a62,
32'h3e95c0fa,
32'h3c254beb,
32'h3d962211,
32'hbea1c81e,
32'hbc630b1b,
32'hbe887d89,
32'hbca2dc75,
32'hbd87abde,
32'hbea52df4,
32'hbe0dfc37,
32'h3ea127dd,
32'hbe6c5d78,
32'h3cb95dca,
32'hbe67d55e,
32'hbd349665,
32'h3ddfc46e,
32'hbe192708,
32'h3e81de7e,
32'hbe214bef,
32'h3eeb7455,
32'hbc37254a,
32'hbe7bce55,
32'hbed88f4f,
32'h3e783267,
32'h3ea72822,
32'h3c99d785,
32'hbe517ca8,
32'hbe107cea,
32'hbe82c6e9,
32'h3e245bf0,
32'h3f018799,
32'hbd3e69ec,
32'hbca56d52,
32'hbe6d7811,
32'h3e25a84c,
32'hbe92c471,
32'hbe697763,
32'hbe13f8ae,
32'hbfb307eb,
32'hbd51eb55,
32'hbe531189,
32'h3b8a1362,
32'h3cc13a6e,
32'hbe2bd503,
32'hbebe0d23,
32'h3e70dfe3,
32'hbdbb9d67,
32'h3dfb75ac,
32'hbead07c1,
32'hbe1e669a,
32'hbef6ed82,
32'h3d9a3205,
32'hbe2cca26,
32'h3e1e951b,
32'h3eb655f5,
32'hbeb119df,
32'hbf066541,
32'h3e1783e0,
32'hbcaff3cc,
32'h3d893029,
32'h3e47b836,
32'hbd33aede,
32'hbcb9fcd1,
32'hbe956d25,
32'hbd2a8939,
32'hbe878559,
32'hbd4fb7b4,
32'hbeee4314,
32'hbf1d7eb9,
32'h3e43e522,
32'hbed3f7f7,
32'h3dedd090,
32'h3e5b59ca,
32'hbe91053e,
32'hbe564e03,
32'h3e6ed2f2,
32'h3e396d2b,
32'hbca740c9,
32'hbe2602ad,
32'hbe93e9bc,
32'hbf0389cf,
32'h3e8fc920,
32'h3dbfcc0f,
32'hbd6cde12,
32'h3f1d6f84,
32'hbe9a16ab,
32'hbe6959cc,
32'h3d9c93c6,
32'hbd7a1ba1,
32'hbe922648,
32'h3d5a55f9,
32'hbde17771,
32'h3ccdb20b,
32'hbe1b654d,
32'h3d6e2dc1,
32'hbe97958e,
32'hbe42cb10,
32'hbd7cd249,
32'h3e34cef2,
32'h3cd7ac69,
32'hbf077cd5,
32'hbeb729c7,
32'h3e812028,
32'hbe0d002e,
32'hbcd2fdfa,
32'hbdfef1b7,
32'h3da5211a,
32'hbdafc3d4,
32'hbd811cbc,
32'hbe38db83,
32'hbf030d3f,
32'h3edcb84c,
32'hbdcb69f3,
32'hbe84f442,
32'h3ef08d02,
32'hbe7834cb,
32'hbe3d880b,
32'h3cf7d6dc,
32'hbd7be09c,
32'hbeda2ddf,
32'hbd6876b5,
32'hbdc179a1,
32'hbd9ab753,
32'hbe33aee0,
32'hbd08ff2e,
32'hbe73784f,
32'hbc93bfbd,
32'h3e9ecfd9,
32'h3eacf3dd,
32'h3e25adae,
32'hbe6b97ec,
32'hbe5dbc82,
32'h3e6b2a24,
32'hbd779c9b,
32'h3d3830d0,
32'h3d89289e,
32'h3e0a2349,
32'hbe851a81,
32'hbd72c46b,
32'hbd5e34cc,
32'hbe76588e,
32'hbd909030,
32'h3aa9dcd4,
32'h3cc6ab31,
32'h3eb2d839,
32'h3e780794,
32'h3ee97f1c,
32'hbd30a5a2,
32'h3e24c8d6,
32'hbe64751b,
32'hbe14c0d0,
32'hbd496c45,
32'h3d625b0a,
32'hbe5fcc83,
32'hbcde3e0e,
32'h3e92e3c6,
32'hbe09ea0e,
32'hbc3e4f8b,
32'h3d98e69f,
32'h3e622f65,
32'hbcb1ddb4,
32'hbe2001e7,
32'hbd84903c,
32'hbf2bb988,
32'hbe22a482,
32'h3dd77e3a,
32'h3ed17f2b,
32'h3d9205ba,
32'hbdc70c69,
32'hbe689c4d,
32'hbef90f4e,
32'hbd3d2484,
32'hbe84172d,
32'hbd85d729,
32'h3e01f2d7,
32'h3e97f453,
32'h3e9e1d11,
32'h3e278f62,
32'hbceda818,
32'h3e70f870,
32'hbe043f55,
32'h3c35eda5,
32'hbbcc2570,
32'hbda1f44c,
32'h3d9d3332,
32'h3e99b302,
32'h3d7c1ca7,
32'h3d079eec,
32'hbcb6f8f1,
32'hbd40ac1d,
32'hbde91b4d,
32'hbeacef91,
32'hbcac99fc,
32'hbfe0172a,
32'h3c8f39d1,
32'h3e24a1b9,
32'h3e4f6323,
32'h3e3f67ad,
32'h3d78b4d7,
32'hbe40dcbc,
32'hbef9e799,
32'h3ccf3584,
32'hbf0daca2,
32'hbe7ec08c,
32'h3e07fdc4,
32'h3def8b18,
32'h3f115b12,
32'h3d3120d4,
32'h3da09cda,
32'h3d58a29c,
32'hbf87f834,
32'hbdb905ba,
32'hbd82c429,
32'hbe20f352,
32'hbe9f43f7,
32'h3e1bdc3f,
32'h3cb35be3,
32'hbde292c0,
32'hbd924295,
32'hbe4ae33d,
32'h3dd6a063,
32'hbe81be05,
32'h3c582985,
32'hbfe89e27,
32'hbcb2c0b9,
32'hbdc46d3e,
32'hbe04f381,
32'h3e05cadb,
32'h3e27fc9a,
32'hbdac3b2d,
32'hbdde1a2b,
32'hbe4ade7d,
32'h3e45e974,
32'hbe956953,
32'hbe18e3fd,
32'hbdf145d8,
32'h3f1760af,
32'h3e93676f,
32'h3d333cfb,
32'hbe401c94,
32'hbdf977d3,
32'hbd6d23e2,
32'hbdcffcea,
32'h3d974d2f,
32'hbdfa394c,
32'hbcb2d237,
32'h3d522491,
32'h3d8e7711,
32'h3ddb7dbd,
32'hbbf58095,
32'h3ebb05d2,
32'hbd89308f,
32'hbd864056,
32'hbf3b6d69,
32'hbd099e80,
32'h3d44c56a,
32'h3ea4d398,
32'hbe1d8566,
32'h3a6f7785,
32'hbe3976d9,
32'hbce9a0b7,
32'hbebfba3b,
32'hbdfa7069,
32'hbdb50e1e,
32'h3d540255,
32'hbd0a1d09,
32'h3e9be845,
32'hbe85460b,
32'h3e9cb563,
32'hbcb7129c,
32'hbdadb1ab,
32'hbc3312cd,
32'hbc72cd2b,
32'hbe869127,
32'h3e6af3b1,
32'h3cc57f57,
32'h3e175301,
32'hbec5f33f,
32'h3ea64d91,
32'hbe9b025a,
32'hbc9b28b9,
32'h3e16d29d,
32'h3e32ac66,
32'hbe474842,
32'hbe1d452a,
32'h3dbdf7da,
32'hbe834f6b,
32'h3e9bc751,
32'h3e30842b,
32'hbeb95182,
32'h3e378624,
32'hbe73c926,
32'h3cbaf31b,
32'h3eb8d053,
32'h3eab9f11,
32'h3dad7fca,
32'h3ec09e14,
32'hc02ee412,
32'hbba56db8,
32'hbf2894a4,
32'h3de9df6a,
32'h3d305fce,
32'h3cc4177a,
32'hbeafa6d1,
32'hbeff9481,
32'h3e8746cc,
32'hbccd8483,
32'hbe88bb24,
32'h3e2d1a0c,
32'hbf4e15cf,
32'h3ead2cd6,
32'h3cd8de4f,
32'h3e9126ed,
32'hbf4d68e6,
32'hbe0f4a64,
32'hbf0902f9,
32'h3ddc716e,
32'h3f0a6a06,
32'h3e88a804,
32'hbfa03bc5,
32'hbf465007,
32'hbf9c6f95,
32'hbd808f77,
32'hbe95f6e8,
32'hbe93aeb6,
32'hbd9fb71d,
32'h3e91c366,
32'hc03f1ba3,
32'h3ea36e50,
32'hbfcde5cb,
32'hbf634b3f,
32'h3d99c60b,
32'h3dae42c7,
32'hbfc1275c,
32'hbf79e1bf,
32'hbfb2b7ed,
32'hbe90f4d3,
32'hbf485fd3,
32'hbf0713ab,
32'hbfab3bf0,
32'h3eeff3a2,
32'h3eb742f9,
32'hbc1eab1f,
32'hbf525909,
32'hbe6b4c5e,
32'hbfa9ca15,
32'h3e6b0e6b,
32'h3f282fa8,
32'h3f3c6d75,
32'hbfa9f312,
32'hbf64be10,
32'hbfd40aa3,
32'hbec031ad,
32'hbf62bb21,
32'hbfdcee8a,
32'h3f2d555b,
32'h3ea5081b,
32'hbfd695c0,
32'h3eaf2bf8,
32'hbf6b39c8,
32'hbf32f882,
32'hbddd10a6,
32'hbd50bccb,
32'hbfcd0165,
32'h3e9c980b,
32'hbf488d43,
32'hbea010a2,
32'hbf9b1575,
32'h3e997dd9,
32'hbfb38d6f,
32'h3e771fed,
32'h3f03bdc5,
32'h3d6afd48,
32'hbef531db,
32'hbe6c7090,
32'hbf8f2784,
32'hbf51abb6,
32'h3eae353f,
32'h3ec7953f,
32'hbe8b29d4,
32'hbf9f9e0f,
32'h3dc3886c,
32'hbf547391,
32'hbe987b14,
32'hbfe3682f,
32'h3eebefb7,
32'h3eadb962,
32'hbf0e3c4c,
32'h3dda82f9,
32'hbdd38d9d,
32'h3ea0abd7,
32'h3c86e31c,
32'hbb9ea319,
32'hbf1d1b51,
32'hbd21ead5,
32'hbf42fac9,
32'h3e11f9cb,
32'h3d54dc4f,
32'hbfc930be,
32'hbee18996,
32'hbe64cde0,
32'hbe8ec988,
32'hbf22a63a,
32'hbe4288ea,
32'hbf26af69,
32'hbf8a8b14,
32'hbf094e0d,
32'h3e9d6d0f,
32'h3e6ef04c,
32'hbc3102cf,
32'hbf8f0f8a,
32'h3e259f77,
32'hbf06d27a,
32'hbe637c8e,
32'hbe99b365,
32'hbd993c4a,
32'h3f22401b,
32'h3e77b71f,
32'hbf3434ec,
32'hbd7b674f,
32'h3db788bf,
32'h3a923564,
32'hbb64b56c,
32'hbe2482f5,
32'hbc643ca0,
32'hbdb91a2f,
32'h3f5642aa,
32'h3d44b8b7,
32'hbf6f1b96,
32'hbf20d0d4,
32'hbf67d90d,
32'hbef143de,
32'hbf6394bf,
32'hbd92978a,
32'hbeb7cd8e,
32'hbd96a9fd,
32'hbebed62f,
32'h3cf20eef,
32'h3e86540d,
32'h3dcdbed7,
32'h3d9dba61,
32'h3c93dfc5,
32'h3d9744a2,
32'hbd0b8153,
32'h3d6f9911,
32'h3db380a5,
32'hbd4514b9,
32'h3dcb9efb,
32'hbc9bde71,
32'h3d7a157e,
32'h3a18d24a,
32'hbcd2a385,
32'hbd793340,
32'h3dbfe82e,
32'hbce3fbce,
32'hbc41b02f,
32'hbe2ddc11,
32'h3c03663a,
32'hbc88e50d,
32'h3e0e9511,
32'h3da1c91f,
32'hbdfde471,
32'hbda4ab18,
32'h3d4e20e1,
32'hbd7f4417,
32'h3b2f7b30,
32'h3d393d48,
32'hbd7cd204,
32'h3e1988bf,
32'h3c45166e,
32'hbdf0211e,
32'h3d2d64ee,
32'h3fb9af82,
32'h3eea2d71,
32'h3d6c3cf8,
32'h3e01a5bc,
32'h3d31469e,
32'h3f4999bf,
32'h3f660b75,
32'hbe8be8a7,
32'h3d8c919d,
32'h3d7ddfc5,
32'h3db7fec9,
32'hbd11c1d8,
32'hbd8a66ad,
32'hbe04ffd2,
32'h3d7994b5,
32'h3d584879,
32'hbe5ea81a,
32'h3f407854,
32'h3e6b7806,
32'hbf9b9625,
32'h3e9acd0b,
32'hbc2d43ff,
32'hbf9c6a41,
32'hbe5dbb01,
32'h3f7f805e,
32'hbdd4243b,
32'h3f24ae69,
32'h3b00ef2f,
32'hbfc24b5f,
32'h3f110c8a,
32'hbf043d95,
32'h3e87488d,
32'h3ec207c5,
32'h3d3057fa,
32'h3ba6b24f,
32'hbf0565f2,
32'hbf0aeb62,
32'hbef8d4aa,
32'h3e35e148,
32'hbda986a9,
32'hbb32de94,
32'h3ea4b490,
32'hbf8e457b,
32'h3d847a97,
32'hbf37dd15,
32'hbea40f84,
32'h3d611b75,
32'h3cad962e,
32'h3eeadbe3,
32'h3ec6f911,
32'h3f399541,
32'h3d96c01c,
32'h3f06fa55,
32'h3cf27040,
32'h3df37dfa,
32'hbe6c72ae,
32'hbc22af09,
32'hbe990067,
32'h3b5b1d7f,
32'h3f42237b,
32'hbd9fd571,
32'hbe95b41b,
32'hbf7e3fcc,
32'h3ee4bbbe,
32'hbee2de79,
32'h3f1c7398,
32'h3e968f26,
32'h3eb115b4,
32'hbf17eb9e,
32'h3c0c07c7,
32'h3be6be71,
32'h3f15486b,
32'hbe672db9,
32'h3e95922a,
32'hbed73c20,
32'h3f6c9b2c,
32'hbe2deff5,
32'h3e75309d,
32'hbe682257,
32'hbf9be4e5,
32'h3e934ab6,
32'h3e21b866,
32'hbd0b802c,
32'h3f279e4b,
32'h3ec1be33,
32'h3edaf4a3,
32'h3d80e533,
32'hbdb0543b,
32'hbfa4e96f,
32'h3eef0b5c,
32'h3e92cea4,
32'h3dceacf3,
32'hbd00d749,
32'hbf5b4eed,
32'hbf4c76ff,
32'h3f349dd0,
32'hbe28ccf2,
32'hbf057f68,
32'hbdbc3baa,
32'hbd18002c,
32'h3d1e9c0c,
32'hbefcee12,
32'h3f132d34,
32'h3e1ba185,
32'hbe45acbc,
32'h3e596f9b,
32'hbe33aad2,
32'h3e6c5632,
32'hbed07da2,
32'hbe388536,
32'hbde22e63,
32'hbc60e4af,
32'h3d5d2439,
32'h3e39ce14,
32'h3ea72f3d,
32'hbe553972,
32'h3d9159ec,
32'hbefd5022,
32'hbf150bc6,
32'h3e7fd64e,
32'h3ebfba18,
32'h3ec19112,
32'hbe3e15ee,
32'hbe457fa6,
32'hbe01ffad,
32'h3f22b6b2,
32'hbd9fec50,
32'h3e347f04,
32'h3e5c46ce,
32'hbd99c16e,
32'hbce32255,
32'hbec0738d,
32'hbe5406d7,
32'hbec6b915,
32'h3e456fa8,
32'hbe5a8aff,
32'h3ed0d7ad,
32'hbe58b3d7,
32'hbc907aeb,
32'hbf2fd550,
32'hbddca024,
32'hbf26aa66,
32'hbd4e3267,
32'hbd3f4fec,
32'hbda24e0f,
32'hbdf2c506,
32'hbf42ba32,
32'h3dcd9617,
32'h3e01f1fc,
32'h3f174f2c,
32'h3e86e5ac,
32'h3c16c01f,
32'hbd3074b7,
32'h3c76979e,
32'h3efad6de,
32'h3e5561d0,
32'h3e97b317,
32'hbe709bed,
32'h3ee39336,
32'hbd8bc41a,
32'hbb94af3f,
32'h3b9427ef,
32'hbf2a82fe,
32'hbcfa28f6,
32'h3e2034b0,
32'hbeef2b38,
32'hbe36050b,
32'h3ecb4c87,
32'hbe314e6e,
32'hbe9d9cc6,
32'h3ea8d6c2,
32'hbf4d71d1,
32'h3d4cab9a,
32'h3d294a1c,
32'h3f0afc2d,
32'h3d96b7ad,
32'hbe485d6a,
32'h3e268323,
32'h3e509443,
32'h3f13fde8,
32'h3e913483,
32'hbded453a,
32'hbe8b696a,
32'h3eae563b,
32'hbedfb487,
32'hbc1308a5,
32'hbef84484,
32'h3d57420b,
32'h3e22815a,
32'h3c8687b2,
32'hbddd807a,
32'hbe092578,
32'hbe9d2899,
32'h3de3e168,
32'h3deb7378,
32'h3e030bda,
32'hbdcf00eb,
32'h3e0277a6,
32'hbe72b2cd,
32'h3e0d8d83,
32'h3ddf0ec0,
32'h3ded483a,
32'h3dbdd708,
32'h3e8daf8e,
32'h3f0c2786,
32'h3d79335d,
32'hbe9ba7de,
32'hbd3e0635,
32'hbe791ace,
32'h3eacc2dd,
32'h3d2632d3,
32'hbdce231b,
32'hbecf9dfb,
32'h3d08658f,
32'hbecbd27e,
32'h3d831b51,
32'hbf41c987,
32'h3dd4161d,
32'hbb8f28e0,
32'hbc9213c6,
32'h3ceb8fb0,
32'hbd281e50,
32'hbe939549,
32'h3e7d6740,
32'h3e31ebfb,
32'hbdcfbd9a,
32'h3e809c4b,
32'hbe08afc6,
32'hbcf3217f,
32'h3c5baee0,
32'h3eca714c,
32'h3e8744ca,
32'hbd5d272c,
32'h3e821058,
32'h3d1acf54,
32'h3d3ff048,
32'hbd32d27a,
32'h3e4bf883,
32'hbdbb172c,
32'h3eca62f6,
32'h3dfcc12d,
32'h3e81b5f8,
32'hbe13ce66,
32'hbdbfb122,
32'h3e14c398,
32'hbef63120,
32'hbf67fecd,
32'h3e5c3180,
32'hbe32fb9a,
32'hbda142f5,
32'hbdb7a827,
32'hbe7fee10,
32'hbdcf4490,
32'hbeab0462,
32'h3e03a135,
32'h3d504f3c,
32'h3d903b04,
32'h3cdc959f,
32'h3dc113c2,
32'hbee2fb2c,
32'h3d1d9c76,
32'hbea66b1e,
32'hbe205a64,
32'h3e415381,
32'h3ed39d59,
32'h3d494851,
32'hbe168fbb,
32'hbc98c1fd,
32'hbd984665,
32'h3ef35c75,
32'hbe961d39,
32'h3e81d43d,
32'h3b958452,
32'hbda59db7,
32'hbdb115c5,
32'hbf800a6a,
32'hbf16366c,
32'h3d08f9fb,
32'hbe282b72,
32'hbdffd976,
32'hbdef8760,
32'hbe48a973,
32'hbec2d396,
32'hbea0ce3c,
32'h3e58bdf9,
32'hbeca2285,
32'hbd1dae0e,
32'h3d8cf83c,
32'hbe67009e,
32'hbda71af6,
32'h3e269c9a,
32'h3cee332c,
32'h3de8e78b,
32'h3d9113ad,
32'h3e81852b,
32'h3de1720c,
32'hbe076b50,
32'hbd15890d,
32'hbf1bd4e0,
32'hbeceef1d,
32'h3d931728,
32'h3e6799a1,
32'hbea22078,
32'hbdee5a02,
32'h3e873cf1,
32'hbf4b8308,
32'hbe937dfa,
32'h3e493bf3,
32'hbec58dd8,
32'h3cecbb15,
32'h38ce2fdb,
32'hbea07dfd,
32'h3e8b3828,
32'hbe2aa6b4,
32'hbd14f55b,
32'hbe9409fe,
32'h3ea3222f,
32'h3c93e769,
32'hbedfab14,
32'hbdd0d714,
32'h3d9b01bd,
32'hbf1c6927,
32'hbcb1998b,
32'h3ecfb477,
32'h3e82b76f,
32'h3e13c65e,
32'h3c4d8fd3,
32'h3e66c33e,
32'hbed897a5,
32'hbef902e4,
32'h3d4f62a6,
32'h3eb5a918,
32'hbde1ec58,
32'hbda8b7cb,
32'hbcd4fd9c,
32'hbf3cfb02,
32'hbed34a5f,
32'h3e17e313,
32'hbdbc1eb7,
32'hbd6ebf14,
32'h3cf4592b,
32'hbe1973dd,
32'h3cdb49ae,
32'hbdbc1a04,
32'h3e183f75,
32'hbc8b85a3,
32'h3e90c6a5,
32'h3e8a7106,
32'hbe322815,
32'hbe901d93,
32'h3e8b8b3f,
32'hbdf248df,
32'h3e25ed89,
32'h3e9d0084,
32'h3ef02441,
32'hbdbc4e51,
32'h3e641437,
32'h3ecc5a81,
32'hbeb22ff5,
32'hbf61cce9,
32'hbde0ae7b,
32'h3c9a8069,
32'h3e43f49f,
32'hbe22f505,
32'h3de7b990,
32'hbe730341,
32'hbde6485f,
32'h3e32a5dc,
32'h3ec31df8,
32'hbd84a599,
32'h3c1d0383,
32'hbdc0f06d,
32'hbea0b608,
32'hbd93b8d7,
32'hbd2f4e91,
32'hbe174a4b,
32'h3db21c8f,
32'hbbbe03d2,
32'h3dfeb840,
32'h3b409b38,
32'h3c1a5fb9,
32'hbdbf4655,
32'h3d8b1dc1,
32'hbe3d5f14,
32'h3ee8b62e,
32'hbe9a89e3,
32'h3e226fd3,
32'h3c87c916,
32'hbe7e018f,
32'hbe93580a,
32'hbd2ee4d9,
32'hbe831a84,
32'h3b8c2fd2,
32'hbc78dd3c,
32'hbde988f4,
32'h3c5c1766,
32'hbdfae22e,
32'h3f09abfa,
32'h3f329e9e,
32'h3d47e63a,
32'hbdbf2ec0,
32'hbde1321f,
32'hbe31d439,
32'hbd9808b8,
32'hbdf50580,
32'hbbf6cefe,
32'hbffd1350,
32'h3e6fbf14,
32'hbf29524f,
32'hbe0a8449,
32'h3e5e6433,
32'h3d24c265,
32'hbd8b160f,
32'hbe50b970,
32'h3e4eac07,
32'hbe2a4a0a,
32'h3aa1a81a,
32'hbd9b497d,
32'hbeab4d45,
32'h3e46465d,
32'hbe3d3dea,
32'hbe5ac154,
32'h3da83a3e,
32'hbd845157,
32'hbf3aad57,
32'h3ecd8497,
32'hbd83ea6e,
32'h3e6a3f6a,
32'h3ea7b257,
32'h3d26f983,
32'hbda5ef48,
32'hbdef67cf,
32'hbe33c17f,
32'hbe8a7acf,
32'hbb897ab4,
32'h3d700a3f,
32'hbdef867f,
32'h3e66cf19,
32'hbf03a596,
32'h3e2a845c,
32'h3eef3c89,
32'hbebd3f78,
32'hbda2661d,
32'h3d066012,
32'h3e4462ac,
32'hbe288fe3,
32'h3e7df715,
32'hbd9524da,
32'h3e199c7a,
32'h3f24db7a,
32'hbe1cb15b,
32'h3d0f8754,
32'h3da63135,
32'h3c990e9d,
32'hbf3b5e11,
32'h3e94f7bd,
32'h3de620e5,
32'hbe040244,
32'h3dc5796b,
32'hbccaeb59,
32'h3cef656d,
32'h3e350fcf,
32'h3dc368d0,
32'hbe8c85d6,
32'h3e3ed82c,
32'h3f02b0a0,
32'h3ef97b86,
32'hbd9cf1f0,
32'hbdb37133,
32'hbe108059,
32'h3df2b743,
32'hbd9a1b22,
32'hbe05ada2,
32'h3d5ddfb4,
32'h3e0b3e10,
32'hbeb06b2f,
32'h3dff7348,
32'hbde06651,
32'hbd8a2ead,
32'h3dd56d8b,
32'h3dc2758e,
32'h3e5aeedd,
32'h3dca3292,
32'h3e3c4641,
32'hbefe2e88,
32'h3e67256e,
32'hbd92dbbd,
32'hbeb0cd9b,
32'hbec45fde,
32'hbd880989,
32'h3d348277,
32'h3d91f9a8,
32'hbd8eaa3b,
32'h3d153434,
32'h3e249134,
32'hbe1bacf0,
32'h3dec86e1,
32'h3e86d4e9,
32'hbddc4a95,
32'h3b2a555a,
32'h3e95dc64,
32'hbef4884c,
32'hbe2ba737,
32'h3e494cfa,
32'h3ed45c0b,
32'hbe7e118b,
32'h3e8bd7a1,
32'hbeca1d50,
32'hbe713a0c,
32'h3dc81a49,
32'h3d4d313a,
32'hbe053e63,
32'h3e8111ee,
32'h3c9cf23f,
32'hbe02c18b,
32'h3e4154cb,
32'h3d044e3a,
32'hbe5c7a5e,
32'hbe4bdc15,
32'hbc0ac062,
32'hbd02bfab,
32'hbe82dd04,
32'h3e4ba039,
32'h3deb2e46,
32'h3e42787a,
32'hbc91738c,
32'hbe007f6a,
32'hbdb0be30,
32'h3d9b7441,
32'hbe66d9b7,
32'h3d34b0d5,
32'hbfe9b47b,
32'hbe015fd7,
32'h3d74f097,
32'h3e386b41,
32'hbe927873,
32'h3ef16a21,
32'hbdc2994f,
32'hbec841d0,
32'hbe0656c6,
32'hbdbfdf50,
32'hbea423c1,
32'h3f17d630,
32'h3e5621e1,
32'h3dd99315,
32'h3e42ebe1,
32'hbdf22db9,
32'hbe4f1545,
32'hbf04ea5e,
32'hbcf01ea2,
32'h3ccc7a41,
32'hbdc22bf8,
32'h3c989c38,
32'h3f0d315d,
32'h3e0c37cd,
32'hbd4643f7,
32'h3c8a53ca,
32'hbd37e8ba,
32'h3c04b069,
32'h3d9bbdd4,
32'hbbc72391,
32'hc0044b40,
32'hbc5f861f,
32'hbe221eb3,
32'h3d45effe,
32'hbe1ec928,
32'h3dc755ef,
32'h3dc2933f,
32'hbeaa6cad,
32'hbec7e5f5,
32'h3bf9d640,
32'hbe40bf78,
32'h3efbca55,
32'h3e0bb652,
32'h3def72e9,
32'h3eb2c7d6,
32'hbd7b08b1,
32'h3e04d249,
32'hbfc280ea,
32'h3cb42ab1,
32'hbcd53f0d,
32'hbd680c57,
32'hbe2dd6ff,
32'h3ea1f87a,
32'hbda465fa,
32'hbf02631e,
32'h3e868840,
32'hbe81aa83,
32'h3eb994a4,
32'h3d3dc1b0,
32'hbe498a50,
32'hbfc42c23,
32'h3d92f9c2,
32'hbceed657,
32'h3e5f2d1e,
32'hbec9a418,
32'h399285e4,
32'hbcb89403,
32'hbe93eb5c,
32'hbdb542a3,
32'h3ec69a71,
32'hbe6fcfea,
32'h3ca4684f,
32'h3d1588fa,
32'h3eb9b866,
32'hbc58d118,
32'hbd2f5626,
32'hbe1e1791,
32'h3eaa7915,
32'h3cea0ae8,
32'hbd69388f,
32'hbe7db265,
32'hbdb3661d,
32'h3ea00c9b,
32'h3e058205,
32'h3d9336bf,
32'h3d742c27,
32'hbe10c799,
32'h3e712d5c,
32'h3e199097,
32'h3d3a4472,
32'hbfb6995b,
32'hbc8e17bc,
32'hbe95b4db,
32'h3eb64a84,
32'hbeee7606,
32'h3e298e2d,
32'hbe737a63,
32'hbf0acf3f,
32'h3e99971c,
32'h3f00b3f7,
32'hbe1bff9b,
32'h3e20387a,
32'hbb97e259,
32'h3f13376d,
32'hbd9cbf32,
32'hbd97f72b,
32'hbe5dd72b,
32'hbedd707f,
32'hbd86ff00,
32'h3cc41078,
32'hbf02e34e,
32'h3d914ebb,
32'hbdd7c68d,
32'h3ea4aa06,
32'h3edc32b4,
32'h3e1f0127,
32'h3d8e64fd,
32'h3e807026,
32'hba077f70,
32'h3d7cd34c,
32'hbf51aaac,
32'hba522869,
32'h3f248662,
32'h3e1d8a27,
32'h3daaec2a,
32'h3f3e2e88,
32'hbef66f24,
32'hbfab1ee0,
32'hbea79a05,
32'h3e821f64,
32'h3e391bbc,
32'h3ee35ce7,
32'hbea06594,
32'h3e746fd0,
32'hbfd6e092,
32'hbe86d3a9,
32'hbd882041,
32'hbe2f1989,
32'h3c908fa5,
32'h3b47df7b,
32'hbe98e3d0,
32'hbe123bdc,
32'h3efed903,
32'hbdeddd4b,
32'hbedbdfa5,
32'hbcb66614,
32'hbe5ca938,
32'h3d29f196,
32'hbd7e109b,
32'hbe26b578,
32'hbf4b4edf,
32'hbe4dd809,
32'h3eb411d6,
32'h3c04e810,
32'h3eba09c0,
32'h3f41f7de,
32'hbf8df9ca,
32'hbfc121d8,
32'hbfe291d5,
32'h3e4e2cf6,
32'hbf138351,
32'hbe90ab69,
32'h3ed02e0f,
32'h3f2f1c13,
32'hc0431bc0,
32'h3ddf22fc,
32'hbe293983,
32'hbee2604c,
32'hbda21590,
32'h3c7caa71,
32'hbf91c095,
32'hbf872e87,
32'h3e62a92a,
32'hbe9303aa,
32'hbefee035,
32'hbf6ef75b,
32'hbe883439,
32'h3ebf0cb7,
32'hbd1e201e,
32'hbd5c4bc2,
32'hbe645f25,
32'hbe9bf0c8,
32'hbff27a7f,
32'hbe7a2f32,
32'h3df04f91,
32'h3f9561a0,
32'hbfb9797d,
32'hbfbba55b,
32'hbfb60a9d,
32'h3d9d7da8,
32'hbf04201f,
32'hc0036eac,
32'h3e2c32b5,
32'h3ed41b33,
32'hbfc37e1c,
32'hbdd0d051,
32'hbe570972,
32'h3c3f089e,
32'hbd56edee,
32'h3cd947a9,
32'hbfc6e4a8,
32'h3ea4da32,
32'hbf63a7e0,
32'hbe58e791,
32'hbe671886,
32'h3f7e9349,
32'hbf85baf9,
32'h3efc8704,
32'hbf59b520,
32'h3f36df09,
32'hbf365a38,
32'hbe63026a,
32'hbf761041,
32'hbf80d034,
32'h3f8f08e1,
32'h3f3b471a,
32'hbf32eaa5,
32'hc00cdfac,
32'h3fa50d23,
32'hbf5f24b5,
32'hbe2223f8,
32'hbfd48781,
32'hbfb45532,
32'h3f861c3b,
32'h3b62a363,
32'h3df905fd,
32'h3ec5a6f7,
32'h3e0b488d,
32'h3d0df296,
32'h3c89d5c7,
32'hbf3b0010,
32'hbf4e32cc,
32'hbe881aaf,
32'h3ea738dd,
32'hbe8f9a89,
32'hbf0073aa,
32'hbda8884d,
32'h3daa48fc,
32'hbf9cdbfe,
32'hbf11bd8d,
32'h3e380a0e,
32'hbe81d729,
32'hbf8470d6,
32'hbe81ec72,
32'h3f4e1c70,
32'h3c0de6c6,
32'h3f2d04b8,
32'hbfccdea3,
32'h3d9dca34,
32'hbed190d9,
32'hbe7481c6,
32'h3dbfc003,
32'hbe9aa0ee,
32'h3f75f7c0,
32'hbd691cfb,
32'h3de506ef,
32'h3eb46027,
32'hbe29d99b,
32'h3c9265de,
32'h3c4fc231,
32'hbf71c29e,
32'h3d58f5d3,
32'hbdc2f4bb,
32'h3f1bb33c,
32'h3c87b5f8,
32'h3e3934dc,
32'hbe3abfd5,
32'hbe73701e,
32'hbf30be27,
32'h3f6b1135,
32'h3d76c62b,
32'hbf7e6857,
32'hbe123a04,
32'hbeb39b1e,
32'h3f8ab666,
32'h3f99a244,
32'h3dd80cc2,
32'hbf8c646a,
32'hbd3b9c72,
32'hbd9be6a4,
32'hbd664a53,
32'h3bd43f72,
32'h3cf16d70,
32'hbdd0911a,
32'hbd1dd7b9,
32'hbd6ba1c6,
32'h3d44e9af,
32'h3d1ae502,
32'hbd925aed,
32'h3da3928a,
32'hbcaacb16,
32'h3d250f56,
32'hbdc4e409,
32'hbdd33fed,
32'h3c4551db,
32'hbca040b1,
32'h3db7987c,
32'h3dbf7ac3,
32'hbd88531d,
32'hb92ed54d,
32'hbd683fd2,
32'hbd935650,
32'hbc0b80d3,
32'h3e06ef16,
32'hbe341795,
32'h3decb070,
32'h3d043eec,
32'hbd220bf8,
32'h3f82bbb0,
32'h3f36c666,
32'h3ed19ac6,
32'hbd1f37fd,
32'hbecfd418,
32'hbcd7c6b0,
32'h3e85a43e,
32'hbe7d94cc,
32'hbe31fe33,
32'h3ef6908c,
32'hbc33e3ac,
32'h3d59b4d6,
32'h3d1b4c3e,
32'h3d55adc0,
32'h3c30eb53,
32'hbe3b9bc6,
32'h3f83a6e4,
32'h3e98bd1a,
32'h3f28003b,
32'h3f0941c5,
32'hbeb57262,
32'hbe36b545,
32'h3dbb0eab,
32'hbf0a9739,
32'hbed7c6fd,
32'h3f03df73,
32'hbf134ad5,
32'h3e247a4c,
32'h3e5bed23,
32'hbf1fc261,
32'h3db13552,
32'hbf027b2b,
32'h3cf694ea,
32'h3e5a3d2c,
32'hbd8dcc94,
32'hbdbee7b8,
32'h3ecb602d,
32'h3e8d0be8,
32'hbefdaa0e,
32'h3e1d15e2,
32'hbce42f7c,
32'hbd5b0fe6,
32'hbe66ef2f,
32'h3e02e8c5,
32'h3d99b745,
32'hbed8c5c3,
32'hbef8f8c5,
32'hbe8645f9,
32'hbe0bd09a,
32'h3eed0457,
32'hbe9d330e,
32'h3f045901,
32'h3da952d3,
32'h3f8d4a82,
32'hbf1c5228,
32'hbe04c95c,
32'h3df28b94,
32'hbb233d75,
32'hbdd7aa4c,
32'hbe02e9a8,
32'h3eb293bc,
32'hbcbaffe4,
32'hbe36d484,
32'hbfbe25a6,
32'h3e34de2d,
32'hbed0fe3b,
32'h3f0f2c99,
32'hbd82d81f,
32'hbbe3f8f5,
32'hbf80fc2a,
32'hbcf31b99,
32'hbd505e0b,
32'h3e290fe1,
32'h3e18ab90,
32'h3e629b09,
32'hbda746b0,
32'h3e8cccd6,
32'h3f10398b,
32'hbda6d48f,
32'h3e535f78,
32'hbeab93bf,
32'h3f216cd0,
32'h3e7f0878,
32'h3e33dab5,
32'h3f4cc0c4,
32'hbf0564b0,
32'h3e769879,
32'h3c0be39c,
32'hbeb149e8,
32'hbeaec1d5,
32'h3f7daf45,
32'h3e2962d0,
32'h3da53401,
32'hbf05a9d0,
32'hbf263686,
32'hbf220fa7,
32'hbec707cf,
32'hbe994b86,
32'hbf2736cf,
32'hbe49d829,
32'hbd529790,
32'hbd006b0e,
32'h3db83331,
32'h3e8895e2,
32'hbd104d58,
32'hbdad0031,
32'h3f59742d,
32'h3d090919,
32'h3eaa596d,
32'hbecc5305,
32'hbef0b227,
32'h3ef0c7ec,
32'h3dc8ae25,
32'h3dcfbe5d,
32'h3ebd38e0,
32'h3f275f89,
32'h3e82fae6,
32'hbec5de2b,
32'hbf2366be,
32'hbed7ec12,
32'h3f1e2046,
32'h3eb60941,
32'h3e54754e,
32'h3b8bb333,
32'h3e688ffe,
32'hbd50412f,
32'hbf86474c,
32'hbd48fa43,
32'h3f89d07b,
32'h3e0bd803,
32'h3dc30099,
32'hbc50d9b5,
32'h3e5ae26a,
32'h3f0a11e2,
32'h3e2480e5,
32'hbb89b928,
32'h3ee376fc,
32'h3dc79a1d,
32'h3c6bd2a6,
32'hbd3a6c07,
32'hbf5b3856,
32'hbd964ec4,
32'hbf7bdc3e,
32'hbef610d8,
32'h3ebff0e4,
32'h3ec8ed56,
32'h3d1f6980,
32'hbd0fddf6,
32'h3e38543f,
32'hbefece4b,
32'h3ed120ff,
32'h3d9db0d6,
32'h3c9f4bc1,
32'hbe475a2a,
32'h3e163fa6,
32'hbeeb95b2,
32'hbf3b00f6,
32'h3eae4abe,
32'h3e589e4c,
32'hbe4a0de3,
32'hbdfcca83,
32'h3db00059,
32'h3ed67a73,
32'hbf38a1f9,
32'hbeaf5e11,
32'h3e4552e2,
32'hbecf7197,
32'hbf26cee2,
32'hbe0dfc67,
32'h3da5f8f2,
32'hbf183f6c,
32'h3eb1fc58,
32'hbf82733e,
32'h3e6aa93e,
32'h3f033604,
32'h3ec57abb,
32'h3e5c26f6,
32'hbdb19690,
32'hbeb9acb8,
32'h3d026c47,
32'h3e08ca4c,
32'h3ccd9330,
32'hbe65d1a5,
32'hbe9e02d9,
32'hbe42d39e,
32'h3e3035e0,
32'hbf8b6fb5,
32'hbeaec4b4,
32'h3e5eaa98,
32'h3daf324e,
32'hbd2825c3,
32'hbdbdb9f5,
32'hbd10d052,
32'hbf002eae,
32'h3e2ecd50,
32'h3e93b312,
32'hbe450d19,
32'h3b3996ac,
32'h3cc19ccf,
32'hbe91284a,
32'h3d2cb58e,
32'h3e84bdac,
32'hbe02551f,
32'h3e8adaae,
32'h3ebe0bf0,
32'h3ab814ec,
32'h3d5e2dfe,
32'hbe859ebd,
32'hbf2dd602,
32'hbed3df21,
32'h3d6b0bf0,
32'hbd86ef23,
32'h3e1a25e5,
32'hbe9a8f1c,
32'hbe0e2f81,
32'hbc99ad8c,
32'hbffcb9e9,
32'hbeddab59,
32'h3df5128e,
32'hbe8ee935,
32'hbd795bc0,
32'h3d2946f3,
32'hbe9f8bea,
32'h3e188312,
32'h3e64d36e,
32'h3c560329,
32'hbe71925e,
32'h3d361b85,
32'h3d9b6306,
32'hbd19a294,
32'h3e3b0e83,
32'h3e3fcbf8,
32'hbf0e8880,
32'hbd1cea84,
32'h3f5984b6,
32'hb9f4d533,
32'h3d8f8f40,
32'h3e13eaf3,
32'hbf61aae7,
32'hbeb89b0f,
32'hbe0e3c24,
32'hbc57251d,
32'h3c30df54,
32'hbdd7a977,
32'hbe020899,
32'h3cfda349,
32'hbff1c497,
32'h3e8ca944,
32'h3e99c011,
32'hbebaf371,
32'hbe00ede9,
32'hbd9dc44f,
32'hbe67e4b7,
32'h3e64397a,
32'hbdbea461,
32'hbde214d5,
32'h3d35f5b2,
32'hbd1c2ea6,
32'h3e58f41d,
32'hbe04f01e,
32'hbe42c7ea,
32'h3e2ec4b0,
32'hbe68f11c,
32'h3c10c794,
32'h3ef2f0b8,
32'h3eb30bee,
32'h3e20bece,
32'hbda0745d,
32'hbf2d8775,
32'hbefe83a7,
32'hbea342f8,
32'h3ca81b6c,
32'hbd2a5c0d,
32'hbeb8fc65,
32'h3c055f8e,
32'h3cb79e9b,
32'hbf8a232c,
32'h3eb77ac4,
32'h3e6bb948,
32'hbc05c106,
32'hbc5c3fa8,
32'h3b993976,
32'hbebe777d,
32'hbe9be1b3,
32'hbe0febcf,
32'h3df9776e,
32'hbf16b11b,
32'h3c032e6e,
32'hbe12222d,
32'hbd9af3a5,
32'h3d5e1e6d,
32'h3da1c18d,
32'hbe84e03c,
32'hbd03340a,
32'h3edbfcb0,
32'h3e31b7b4,
32'h3cb180cb,
32'h3e4e8d43,
32'hbead9cd1,
32'hbf285d83,
32'hbf0c6742,
32'h3f3d4483,
32'hbe076349,
32'hbe8c42f2,
32'hbe28ea42,
32'h3df73971,
32'hbf289f8c,
32'h3d59fa3d,
32'h3ea039ce,
32'hbe5cd9d4,
32'hbb692922,
32'h3d05205b,
32'hbeb47225,
32'hbedbc1f4,
32'h3e0fd5bc,
32'hbd532a09,
32'hbf7e0902,
32'hbb1aeb5c,
32'h3dbc1905,
32'hbe124f35,
32'hbe15984e,
32'h3d524e87,
32'hbda8a41e,
32'hbdf51649,
32'hbe5d36d4,
32'h3e602d9b,
32'hbe3c962b,
32'h3e89c65a,
32'hbeb19851,
32'hbe20a359,
32'hbecf1c64,
32'h3e39d253,
32'hbd67ae38,
32'h3db68c21,
32'hbe6090cb,
32'hbc2180f3,
32'hbeb487f4,
32'hbdc3041c,
32'h3e143828,
32'hbee0cf06,
32'hbd9a6e73,
32'h3c4eb1df,
32'hbf1807e6,
32'hbe097374,
32'h3ec812e7,
32'h3e56ad36,
32'hbe2ac5c3,
32'h3eccc7c7,
32'h3d66a23f,
32'h3e2fcab9,
32'hbd377a7c,
32'h3e7cb7ff,
32'hbe811458,
32'h3e7dbf9c,
32'hbf0fc2eb,
32'h3d5ae20d,
32'hbd3a6f7c,
32'h3d875302,
32'hbe871293,
32'hbc8f49d4,
32'hbf3dc61a,
32'h3dca6b6f,
32'hbec86d05,
32'hbe8e37ed,
32'hbd914523,
32'h3e99c41c,
32'h3ee7d415,
32'h3e86a98f,
32'hbe1dff5c,
32'h3f3e517b,
32'hbcf756f1,
32'hbc0a7aa7,
32'hbe8437fd,
32'hbf49e1e4,
32'h3ec506c2,
32'hbe20f532,
32'hbe88fa1c,
32'hbf26303b,
32'hbdc5d2c3,
32'h3dc1af0c,
32'hbe10f76b,
32'h3e47b5bf,
32'hbe2829d9,
32'h3daf9f6e,
32'hbfa31146,
32'h3cda4cda,
32'hbe9e41ea,
32'h3ea2b2a6,
32'hbf1722ec,
32'hbdb0c23f,
32'hbe1cf331,
32'hbe1ddbe3,
32'hbf5a00ad,
32'h3ec8b47c,
32'hbf2832b2,
32'h3bb6631e,
32'h3f0097a0,
32'h3db6dfa6,
32'h3e49db3f,
32'h3f1b88ad,
32'hbcfa7662,
32'h3d3bd644,
32'hbd6956bd,
32'hbeea169c,
32'hbea6c663,
32'h3e30a353,
32'h3ea4f1ae,
32'hbff7c1f8,
32'hbd468c10,
32'hbf2365b3,
32'hbe230d27,
32'h3e9b7456,
32'hbea86771,
32'h3e3147e1,
32'hbf629781,
32'hbefb064e,
32'hbeaf496a,
32'h3d7a56af,
32'h3cfe9447,
32'hbdfbea48,
32'h3ec10ffe,
32'hbdd4ad84,
32'hbed12fb2,
32'h3e8844b4,
32'hbea0f4f1,
32'hbeaad13d,
32'h3e5c7ead,
32'h3b027eaa,
32'h3e97e122,
32'h3ef1a471,
32'hbe13e5be,
32'hbdcc6a07,
32'h3d32c948,
32'hbf2c2ff9,
32'hbf24db9e,
32'h3dd64299,
32'h3d8bcaa7,
32'hbe3ade14,
32'h3d8ee73b,
32'hbf5a2793,
32'h3e8eb355,
32'h3c9ce46d,
32'hbe97dab6,
32'h3d233874,
32'hbd972e80,
32'h3dc2307f,
32'hbef58123,
32'h3e193168,
32'h3e8915b3,
32'h3e0d04bb,
32'h3f17b11f,
32'hbe09b1f9,
32'hbbab0bc4,
32'hbd5b6595,
32'hbe46f51b,
32'hbf6e3d5b,
32'h3e10a632,
32'h3d88148f,
32'h3eb62943,
32'h3d2ed93b,
32'hbd2b8cf8,
32'hbda31057,
32'h3e08d4e0,
32'hbdce96ce,
32'hbef5d56b,
32'h3e9d7db7,
32'h3e7618f8,
32'h3ded92f7,
32'h3ea08e67,
32'hbdd43e79,
32'hbe1fd8a6,
32'hbc00ce53,
32'hbf92cc48,
32'hbd029a98,
32'h3b9d2d20,
32'h3e8a8e44,
32'hbef0e7af,
32'h3e4d0ae0,
32'h3d8d7f78,
32'h3db63880,
32'h3ec0e682,
32'hbe094e25,
32'h3d54f4c3,
32'h3e24cf91,
32'h3e92cebd,
32'hbf9dcfae,
32'hbba284d9,
32'hbdf91225,
32'h3e1fbe18,
32'hbdd4f9c3,
32'h3c596a95,
32'h3cad302b,
32'h3eea9bef,
32'hbdc74173,
32'hbd2a11a0,
32'h3ee4cc55,
32'h3e900eec,
32'h3e7c2ef7,
32'h3d7ad36f,
32'h3ef398aa,
32'h3bb75971,
32'h3c84db39,
32'hbf9b4de6,
32'h3e2489e4,
32'hbce0df39,
32'h3e94c20e,
32'hbf0596b5,
32'h3e8083ef,
32'h3d8a0741,
32'hbd68042c,
32'h3e27fd73,
32'h3e0f8f39,
32'h3e059280,
32'h3e89ef90,
32'h3dae7cea,
32'hc00c0efd,
32'h3d41b3da,
32'hbe8ad238,
32'hbca38f92,
32'hbea2230b,
32'h3c098355,
32'hbca5bdc9,
32'hbd1429cb,
32'hbb9b79b8,
32'h3e039dac,
32'h3ed84022,
32'h3dbee919,
32'hbc1bd7bc,
32'h3ce282a7,
32'h3e6920bc,
32'h3d77dd54,
32'hbda977fd,
32'hbfc5d1f6,
32'h3d19a44f,
32'h3e15e3ef,
32'h3def4e9e,
32'hbe7beda0,
32'h3e8f76cd,
32'h3e2b3f6a,
32'hbe890526,
32'hbddbd597,
32'h3e539a4b,
32'hbe35d447,
32'h3e15713e,
32'h3e93b4e7,
32'hbfd08d1b,
32'h3e292959,
32'h3dfc2bd0,
32'hbe52fd81,
32'hbf92bd13,
32'hbe2e0546,
32'h3c9207a7,
32'hbd7b618c,
32'hbdc7cebe,
32'h3e02cd73,
32'h3ef1975a,
32'hbd9fafe2,
32'h3e28990d,
32'hbcec803a,
32'h3e2a3c6e,
32'hbd0d1bbf,
32'hbd89db40,
32'hbfb7a48e,
32'hbc606000,
32'h3cc258f1,
32'h3e640b61,
32'hbe9520d2,
32'h3edb6dd3,
32'h3e7db5fb,
32'hbebcbd41,
32'hbee1e3d8,
32'h3dabf581,
32'hbd9c0968,
32'h3e549e1a,
32'hbc91fd84,
32'hbf1408d5,
32'hbe2308a9,
32'hbd9456df,
32'hbed985bb,
32'hbf7d0aec,
32'hbd97213b,
32'h3b8f2d7e,
32'h3d909a3f,
32'hbe83331d,
32'h3e87ecd0,
32'h3e5c5ecc,
32'hbe580f43,
32'hbe259fdc,
32'hbd50518f,
32'h3e5a3139,
32'h3e037b45,
32'hbe5b091a,
32'hbe5220a6,
32'h3c775032,
32'h3e8a495e,
32'h3e200757,
32'hbef12864,
32'h3ed3378e,
32'h3e185723,
32'hbebd43ce,
32'h3ed77ccd,
32'h3e7626c2,
32'hbe98a3fb,
32'h3e9c5403,
32'hbe39b1ef,
32'hbf184cd5,
32'hbebedb25,
32'h3e58cbe2,
32'h3d1089fb,
32'hbe855cce,
32'h3add375e,
32'hbcb4b75a,
32'hbd3439e6,
32'hbe014f77,
32'h3ec0a0c8,
32'h3da217f8,
32'h3e44ecf1,
32'hbe5fd773,
32'hbe84ced5,
32'h3df77db6,
32'hbe027d44,
32'hbd756245,
32'hbfbcbcdb,
32'hbd27ccc3,
32'h3e837599,
32'h3d976e8f,
32'hbea34e48,
32'h3f170653,
32'hbd55e0d1,
32'hbf1d88dd,
32'h3e179664,
32'h3ec3cec0,
32'hbe549155,
32'h3f0d151f,
32'hbe457468,
32'hbe9015cb,
32'hbe89b51f,
32'h3e542799,
32'h3d5c0856,
32'h3f6bcf27,
32'hbc88edda,
32'hbd4d3c17,
32'hbe65c6c2,
32'hbd77bd63,
32'hbe971f7f,
32'h3ee74a31,
32'hbef37772,
32'hbe33e29b,
32'hbc742a05,
32'hbe63ddf7,
32'hbd512e88,
32'hbe8a8d5e,
32'hbf95c04c,
32'hbe04237d,
32'hbe58f3bd,
32'h3d7a2c62,
32'hbf12e1cb,
32'h3f33e709,
32'hbdcea2e0,
32'hbf28d67a,
32'hbf4b1009,
32'h3ef64bb1,
32'hbe0e3e70,
32'h3f43eae6,
32'h3d9a765b,
32'hbf19de3e,
32'hbfc33885,
32'hbe3ab83d,
32'hbe106199,
32'hbe6d4c67,
32'h3d6856b7,
32'hbc9b3d91,
32'hbed8cf87,
32'hbf696d53,
32'h3e2f135f,
32'h3e8416e4,
32'hbf26eb7e,
32'hbf065364,
32'hbed0021c,
32'hbee45bca,
32'hbdd35307,
32'hbdfef19b,
32'hbf647682,
32'h3e6eeccb,
32'hbf261954,
32'hbea563e5,
32'h3e313fc9,
32'h3f4cced6,
32'hbfad2173,
32'hbfa94ecb,
32'hc0176839,
32'hbe90ec51,
32'h3eec7a93,
32'hbd802acc,
32'h3dee0d17,
32'h3d99f8ae,
32'hbfcc1c87,
32'h3ea24fb9,
32'hbebff066,
32'hbf02e128,
32'hbdf40adc,
32'h3987576a,
32'hbf82b69f,
32'hbf2360c3,
32'h3f47c212,
32'hbeb6b889,
32'hbf10e118,
32'h3f002a47,
32'hbecb6eff,
32'h3ec916ba,
32'hbf097e87,
32'h3eb25535,
32'hbf020d02,
32'hbe48247f,
32'hbf19ad98,
32'h3e8af643,
32'h3c9a2fe3,
32'h3f814a75,
32'hbf818369,
32'hbfb19cd3,
32'hbf927d38,
32'h3e9f084b,
32'hbe8d74c3,
32'hbf99ed51,
32'h3e868701,
32'h3e9820e1,
32'hbef74eb4,
32'h3f126118,
32'hbeb13d2b,
32'h3f216651,
32'hbcf4af0c,
32'h3d808050,
32'hbf5e34f1,
32'hbe89ceed,
32'hbf078871,
32'hbe12c58c,
32'hbee2c3f9,
32'h3f525419,
32'h3eda73bc,
32'h3da0bfef,
32'h3ed3f54e,
32'h3eaaa905,
32'hbf4a9d07,
32'hbf126617,
32'h3b8344f2,
32'h3c210b57,
32'hbda88a1c,
32'h3f799872,
32'hbf2311df,
32'hbf7dc67a,
32'h3f1bf88e,
32'hbf2a58b6,
32'h3ebdca5a,
32'hbf9ff3af,
32'hbfb043b2,
32'h3f4c8208,
32'h3e1d75b3,
32'hbebb9d0e,
32'hbe66651c,
32'hbd9f1ea7,
32'hbbf3aba8,
32'hbcd82d5c,
32'hbf228c41,
32'h3db79504,
32'h3ec612f6,
32'hbe48866b,
32'hbe8a3a6a,
32'hbecbc545,
32'hbf543d79,
32'hbda8446b,
32'hc0031a92,
32'hbdc2bd06,
32'h3e319023,
32'hbee010e0,
32'h3eca1f30,
32'hbee571c3,
32'h3f694e16,
32'h3ee53534,
32'h3ea280ee,
32'hbfa4f1e8,
32'h3f315c20,
32'hbef033ba,
32'hbe05c178,
32'hbdadc4fd,
32'h3d465a68,
32'h3f8806f7,
32'hbe0b9cf0,
32'h3d144d4a,
32'h3df21675,
32'h3f1851c6,
32'hbd7e4bcc,
32'hbca3a0f1,
32'hbe5d4642,
32'h3d6d39c0,
32'hbbb503fb,
32'h3e894072,
32'hbc6ba180,
32'h3e2bd66c,
32'hbe431637,
32'hbdad9ad2,
32'hbe58208d,
32'h3e0415c6,
32'hbd3aefe8,
32'hbf191c9d,
32'hbdf5d0ac,
32'hbd4945f5,
32'h3eb05b2a,
32'h3f05f9a5,
32'h3d3601cc,
32'hbedd837d,
32'h3d4ae9b0,
32'hbb8b3d0f,
32'h3d25634b,
32'h3da4c3b5,
32'h3d13bec5,
32'hbb269434,
32'hbdbcddec,
32'hbda55163,
32'h3d594099,
32'hbc510feb,
32'hbca34627,
32'h3da28dd0,
32'h3d6bccf0,
32'hbd1b9b93,
32'hbd53a9b1,
32'hbd97a569,
32'hbd3a1cec,
32'hbcbbbcda,
32'h3e1cd853,
32'h3e455eaa,
32'hbda0e3c0,
32'h3cd234eb,
32'hbd32157c,
32'hbde14537,
32'hbd1f70de,
32'h3d28d4da,
32'hbe1a0276,
32'h3e28c3cf,
32'hbd8d1040,
32'hbdbedf06,
32'h3e27f6fc,
32'h3f433a69,
32'h3e8de4d9,
32'h3ec4ebdb,
32'hbf16e5f5,
32'hbe1fb886,
32'hbd384c58,
32'h3dc6599f,
32'hbe516c32,
32'h3e5976c2,
32'h39a37923,
32'hbcd196c1,
32'h3f468b59,
32'hbded2e4e,
32'hbd7554a8,
32'hbf3d3686,
32'h3e58ffce,
32'hbeb085bc,
32'hbe68b9da,
32'h3d74cba1,
32'hbdd0e697,
32'h3f1269ae,
32'hbccffc45,
32'h3ebc5e93,
32'hbe6908b2,
32'h3f89d9fa,
32'hbe816f44,
32'h3ead1298,
32'h3d12cc61,
32'hbe919f02,
32'h3e1c1bd1,
32'h3ef6c1e2,
32'hbe444124,
32'h3da0c5e2,
32'h3e04fe94,
32'h3e5c84b2,
32'hbed28050,
32'hbd79070e,
32'hbf2a87f4,
32'h3f1a54a6,
32'hbde7f304,
32'hbd1fc9ab,
32'h3ec3c5f7,
32'hbf0aa30e,
32'hbf16b590,
32'hbd7897de,
32'hbe90f964,
32'hbed87b57,
32'h3f0e782f,
32'hbeadcf72,
32'hbf295832,
32'h3dd118fe,
32'h3ce98e84,
32'h3f122e52,
32'hbf8aa8d0,
32'h3f0eb980,
32'hbeecf934,
32'h3ec8aa4d,
32'hbf15918a,
32'hbf066df6,
32'hbe8c7106,
32'h3f5b95e0,
32'h3dd693d2,
32'hbf854779,
32'hbde95d4f,
32'h3f3adea1,
32'hbf732fce,
32'h3e90f8e2,
32'h3e89e368,
32'hbf192b19,
32'hbc79fd12,
32'h3cd70e75,
32'hbf6a1b9b,
32'hbecaaf39,
32'h3dc43478,
32'h3ea476d8,
32'h3e7c93dc,
32'h3ee8c9f8,
32'h3f33f75e,
32'hbe6c65e2,
32'hbf7e3315,
32'hbe18eaa9,
32'hbf5d25eb,
32'hbe5b12ad,
32'h3e3946af,
32'h3e1117bc,
32'h3e1a1244,
32'h3e414400,
32'hbf1fabf8,
32'h3e629d48,
32'h3f2d31c7,
32'h3e10f153,
32'h3f146929,
32'hbdcf6dce,
32'hbed73983,
32'h3f0e5bd8,
32'hbf979bf8,
32'h3e149c6f,
32'hbf573744,
32'hbd5fe356,
32'hbd283d0e,
32'h39eb873f,
32'hbf18622a,
32'hbec3f784,
32'h3dc511a3,
32'hbe671fd9,
32'h3f90e5a9,
32'hbdcd42b8,
32'h3e2cb164,
32'hbe208c47,
32'hbef4b667,
32'h3e375cc4,
32'hbf17314c,
32'h3d667b9f,
32'h3f371f92,
32'h3ee1aa5d,
32'h3f21be04,
32'hbe83dd4d,
32'hbf5df682,
32'hbeaea75c,
32'hbb012161,
32'h3dfa160c,
32'h3e05f6a1,
32'hbf197ee3,
32'hbe4732df,
32'hbe0d610b,
32'hbfe689fb,
32'hbe593ae7,
32'h3ee4fe35,
32'h3ecc199f,
32'h3c9ce0c7,
32'h3bca23c7,
32'hbec32fd4,
32'hbe9a2851,
32'h3de7a879,
32'h3eadf6f7,
32'h3f374268,
32'h3e54019c,
32'h3e5d25c8,
32'h3d2e8b02,
32'hbe31a297,
32'hbdf6234f,
32'hbea9d4c8,
32'hbe6ab0a6,
32'hba9d49f1,
32'h3dab8965,
32'hbde4b481,
32'hbee9cd6d,
32'hbf46507e,
32'h3df00df9,
32'hbe90f8ae,
32'h3c8c5a1e,
32'h3ec8f1f6,
32'hbf0031dd,
32'h3d5fa898,
32'hbcc914eb,
32'hbfc85de8,
32'hbe7568e5,
32'hbd82fef4,
32'h3d10843f,
32'hbd82e888,
32'hbdabf5c8,
32'hbdd2e1f8,
32'hbf6cc677,
32'hbe38670d,
32'h3dcead04,
32'h3f15f99e,
32'h3d9a8cde,
32'h3e0d6d01,
32'h3dda37aa,
32'h3e0a10c0,
32'h3e0ada62,
32'hbecb356b,
32'h3e7b5b09,
32'h3f393a3e,
32'h3e9245df,
32'h3e28a4ad,
32'hbe7f9917,
32'hbf6bd1a6,
32'h3d05131b,
32'hbf28f947,
32'h3d0b3c44,
32'h3e90d5c9,
32'h3d3e085e,
32'hbe16371c,
32'h3ed47b15,
32'hbfcf65f9,
32'h3f040306,
32'h3ee16b6c,
32'hbe1100b0,
32'h3cae69e0,
32'hbd5d545c,
32'hbe514a5c,
32'hbf4b35f3,
32'hbe17a034,
32'h3e51adce,
32'h3e826245,
32'h3b03b0c4,
32'h3e8d42c9,
32'h3c96bfe7,
32'hbe1cac34,
32'hbd68be75,
32'hbf085d01,
32'hbc4cc3ef,
32'h3f19ac41,
32'hbda4d6e7,
32'hbc8d70f2,
32'hbdcf4675,
32'hbfaa95a0,
32'h3e1ee4f8,
32'hbf019c99,
32'hbe6a8cf1,
32'h3ed37bc5,
32'hbd410bbd,
32'hbcc62472,
32'h3ac0af02,
32'hbf9e4ee2,
32'h3f2d5b92,
32'h3ec94a15,
32'hbe974a5d,
32'hbd98be61,
32'hbd7331a8,
32'hbecfc643,
32'hbfa47f81,
32'hbde75b8f,
32'h3e849293,
32'hbeac1719,
32'h3b3b415c,
32'h3e6bf73a,
32'h3e2afa49,
32'h3ec1ee8f,
32'hbd906588,
32'hbeb2b5fb,
32'hbe1d29c5,
32'hbdd497f8,
32'hbd866426,
32'hbd699370,
32'h3d758c99,
32'hbfaf3fd6,
32'h3e740cfc,
32'hbde2e879,
32'h3e75025a,
32'h3e331574,
32'hbe8227e3,
32'h3d7f130d,
32'hbeb8c4ea,
32'hbf2a434c,
32'h3e1af948,
32'h3ed4ff06,
32'hbec7e0a9,
32'hbc162805,
32'h3cc1dbba,
32'hbe8e3163,
32'hbfc2bba9,
32'h3e815cda,
32'h3dfd7729,
32'hbe083a44,
32'h3e4bedef,
32'h3d8e29c7,
32'h3bd61140,
32'h3e090207,
32'h3d73f540,
32'h3e6dca94,
32'hbdb3c4b0,
32'hbfac8007,
32'h3dbd8716,
32'hbd839483,
32'h3d443846,
32'hbf829186,
32'hbb95849b,
32'hbe6e3dbe,
32'h3ec1fb86,
32'h3eb38298,
32'h3d5b9299,
32'h3df8060d,
32'hbd32c8cc,
32'hbe72a7e6,
32'h3e1d1ee1,
32'h3ee3b93c,
32'hbd5e7a93,
32'h3ce7e025,
32'hbd5dab2a,
32'h3e7b5387,
32'hbf949f51,
32'h3efb4405,
32'hbd9d0573,
32'hbec9f579,
32'h3eaf591b,
32'h3de39d04,
32'h3e38a238,
32'h3e7f4ea4,
32'hbd9a4e95,
32'h3d39ec7d,
32'hbc39ba44,
32'hc01b3775,
32'h3e38da53,
32'hbddbbee5,
32'hbaee96d0,
32'hbf8f48cb,
32'h3c6715a7,
32'hbef14417,
32'h3eb28b93,
32'h3ef43bcf,
32'h3de5f433,
32'h3d8924b5,
32'h3d2d9dbd,
32'h3d9fef36,
32'h3e6b387d,
32'h3f231635,
32'hbe3e3047,
32'h3d4121c0,
32'h3cf8da30,
32'hbe536300,
32'hbf51fdd1,
32'h3ee5ca4e,
32'hbd33a9b9,
32'h3e2996bd,
32'h3dd1cd8d,
32'h3de2a4ba,
32'h3e20d16a,
32'hbe13954d,
32'hbd8f96d1,
32'h3dac25b7,
32'h3d22a3b6,
32'hc02c04a4,
32'h3ec0b2ca,
32'h3db2d3de,
32'hbd7b25f9,
32'hbf3f79ce,
32'hbd48ccf9,
32'h3e0a19c1,
32'h3ef81723,
32'hbf341381,
32'hbee2d1fd,
32'h3e287282,
32'h3e631b69,
32'h3f0a2059,
32'h3dc166f7,
32'h3eb8d256,
32'hbddd1ec4,
32'hbde5decb,
32'h3b04c0b7,
32'hbeeee530,
32'hbfa40d79,
32'h3efb1677,
32'hbd28ac4f,
32'hbe1b46c6,
32'h3ea3cbe7,
32'h3b86e8d7,
32'h3ec43c7c,
32'h3e5a1d4b,
32'h3e79fd09,
32'h3e614ae1,
32'h3dbcb2d2,
32'hbfe22465,
32'hbdda27d5,
32'hbd27d51a,
32'h3e23dfce,
32'hbf2042d0,
32'h3e377ad7,
32'hbef4d353,
32'h3d1639c1,
32'hbfa46cf8,
32'hbdd5cd02,
32'h3e30ae8b,
32'h3ea8deb5,
32'h3e9ad78f,
32'h3e916737,
32'h3d9b3739,
32'h3ea0eb0c,
32'hbc485c3f,
32'hbc83d721,
32'hbe0552d7,
32'hbf80f47b,
32'h3c56d486,
32'hbe14a4bc,
32'hbeb076a8,
32'hbf9369ce,
32'hbe10763f,
32'h3e10e68d,
32'hbe884969,
32'h3e14483a,
32'hbd51fe24,
32'h3e887765,
32'hbeb4bb91,
32'hbef45e01,
32'hbd6b277b,
32'h3d4dcc0a,
32'hbece786d,
32'hbe55aa6d,
32'h3e2d02ab,
32'hbd71a5ec,
32'hbf0855d2,
32'hbead4723,
32'hbefa2e93,
32'hbd9d6a6e,
32'h3ebc5c74,
32'h3ec3e100,
32'h3e779912,
32'h3e9ee83c,
32'h3d06301e,
32'hbda3f55c,
32'hbe83599c,
32'hbe458d54,
32'hbebccfb0,
32'h3e4ce532,
32'hbdddc0a5,
32'hbf94dedf,
32'h3e176760,
32'hbf00f97a,
32'hbe6a68d9,
32'h3d46c963,
32'hbe48b1b3,
32'h3d1045b7,
32'hbe02fc22,
32'hbab5ffeb,
32'hbe1768d6,
32'hbbea1209,
32'hbd5f6526,
32'hbdded7d6,
32'h3f240a23,
32'hbedcb435,
32'h3e3895d2,
32'hbf34de8e,
32'hbdf9fe3f,
32'h3e190db9,
32'h3e0cf6d2,
32'h3f1bd359,
32'hbc3f6eec,
32'h3edd7233,
32'hbcef2c35,
32'hbceba427,
32'hbf007f72,
32'hbf172838,
32'hbecaa9be,
32'h3d31b996,
32'h3e398a6b,
32'hbdeafdc2,
32'h3eb5ed02,
32'hbf29409b,
32'h3d075c77,
32'hbda97b03,
32'hbf1111c5,
32'hbe99ae0e,
32'h3e572f0e,
32'h3de9c026,
32'hbddb6550,
32'hbeb66b65,
32'hbd85b681,
32'hbdff423c,
32'h3e64d6aa,
32'hbe532ca9,
32'hbe659b39,
32'hbf7f2394,
32'hbe18584a,
32'hbdc2f782,
32'hbec06dae,
32'h3e6f2b0f,
32'h3d5d56a2,
32'h3e660ee6,
32'hbb52f4a6,
32'hbddfe9ba,
32'h3e170ec0,
32'hbec5847d,
32'hbf1eb679,
32'h3e8380ac,
32'h3e8e6bc2,
32'h3ece9ca0,
32'h3d953df3,
32'h3e800e00,
32'hbc91ae6a,
32'h3eaef1ba,
32'hbf4b1687,
32'h3ea3b21d,
32'h3d9c4773,
32'hbd46157b,
32'hbd8e9e1a,
32'hbf040288,
32'h3e352ab4,
32'h3e568482,
32'h3e5c1c8b,
32'h3cd44e25,
32'hbddda3a5,
32'hbf6cf3ba,
32'h3e956c3f,
32'hbe31bb1c,
32'hbe053443,
32'h3e222894,
32'h3d011000,
32'hbe8f5ed8,
32'hbd81980e,
32'h3c37d876,
32'h3d71997e,
32'hbeb1764b,
32'hbeb90b1c,
32'h3e365859,
32'h3e160740,
32'h3df02d04,
32'h3eab5b14,
32'h3e5ebd57,
32'hbdbae302,
32'h3e94d081,
32'hbf246a37,
32'h3d21e71d,
32'h3b637ba5,
32'h3ebb4279,
32'hbe8c82b1,
32'hbf0492ba,
32'h3e3dc7de,
32'hbc4f683d,
32'h3e862f97,
32'h3e8e1e80,
32'hbdf8c3f6,
32'h3e20b78f,
32'h3e6740e7,
32'hbf6850ba,
32'hbcd2d1fb,
32'h3e3b3f3f,
32'h3d302f75,
32'hbed7d6aa,
32'hbd49d833,
32'hbddc9eeb,
32'hbd7d9454,
32'hbe81b95c,
32'h3e0126b6,
32'h3e87c8b3,
32'h3f00b3e8,
32'hbb222f9a,
32'h3d4892b2,
32'h3eb3b992,
32'hbe63d290,
32'h3d1b89fe,
32'hbe631c51,
32'hbdcb3747,
32'hbd13e7fa,
32'h3df05b59,
32'hbdd2b11d,
32'hbf11bded,
32'h3d918b63,
32'hbe94d798,
32'hbe34311a,
32'h3f10c482,
32'h3e3cad5d,
32'h3ee7c59c,
32'hbe1758ee,
32'hc0106f98,
32'hbde4ccc2,
32'h3e841a33,
32'hbe5965fd,
32'hbed953f0,
32'hbd532f1e,
32'h3a1ad469,
32'h3eacf8e5,
32'hbd09c65b,
32'h3e4a0a6f,
32'h3e433841,
32'hbe83b285,
32'hbdd199ab,
32'h3da7caf1,
32'h3dd6e3fc,
32'hbe9de80a,
32'hbe4a5de2,
32'h3e346c3b,
32'h3e59ddc7,
32'hbe2a0438,
32'h3ea45a89,
32'hbe67c245,
32'hbf069dff,
32'h3e811917,
32'hbf30253b,
32'h3e73d2e2,
32'h3e214367,
32'h3dadee60,
32'h3d90bc58,
32'h3e6371e2,
32'hc00d4a14,
32'hbe63bbc6,
32'h3e5bf337,
32'hbedde59d,
32'hbe58db1e,
32'hbdbe3cb0,
32'hbd89d561,
32'hbe80329c,
32'h3e3242cd,
32'h3cb2a4a7,
32'h3e3812b4,
32'hbe56e1e2,
32'hbe6920a5,
32'h3e0dee8a,
32'h3db39beb,
32'hbe6d5778,
32'hbca52045,
32'hbede2e3a,
32'h3c8135f1,
32'h3ebe32f0,
32'h3eb0907b,
32'hbef87549,
32'hbe1bcfe0,
32'hbcaf6c68,
32'hbf278ca0,
32'h3d5fbe70,
32'hbdeff667,
32'hbec9ca50,
32'h3d967f18,
32'hbcd7f526,
32'hbfdc3bc6,
32'hbf0c6194,
32'h3e3d355e,
32'h3da5b2b3,
32'h3d9dc6ca,
32'h3d6ce099,
32'hbb4d6db6,
32'h3e4e1385,
32'hbe523d47,
32'h3d3f34e7,
32'h3ee84a42,
32'hbee739a7,
32'hbe916d95,
32'h3e8050e1,
32'h3e2f0415,
32'h3e95184a,
32'hbd54d490,
32'hbf14f320,
32'h3eb393ac,
32'h3dd3e58b,
32'hbee42373,
32'hbf0f3ffd,
32'h3e26e032,
32'hbdd1db46,
32'hbe9669ae,
32'hbf593ce8,
32'h3e06f03c,
32'h3e1f1bd1,
32'h3ec423f4,
32'hbd2dff18,
32'hbf938e59,
32'hbf90b87b,
32'h3ce6e801,
32'hbe4624d0,
32'h3eb7ca94,
32'hbddbbfd2,
32'h3d4b0ba7,
32'h3d82dc7a,
32'hbd323305,
32'h3dd777fb,
32'h3f3e38d1,
32'hbfacff73,
32'hbe4544eb,
32'h3e5f6e5b,
32'hbd42fbcd,
32'h3a1883a5,
32'hbe5edf48,
32'hbf056293,
32'h3e88892a,
32'hbf143210,
32'hbf08d313,
32'hbedc71b0,
32'h3f5eeab6,
32'hbe8c7ff0,
32'hbf3d27f0,
32'hbed9f807,
32'h3ece51d0,
32'h3dec6156,
32'h3f106814,
32'h3db83671,
32'hbf29db23,
32'hbf3e742a,
32'h3dea6f58,
32'hbf4f91f6,
32'h3f15aa89,
32'h3d897e30,
32'hbca76121,
32'hbdc7dc52,
32'h3e428755,
32'h3dbe7523,
32'h3e81e556,
32'hbf0e8cd0,
32'hbefc466b,
32'hbe0efb8b,
32'hbe0ccc87,
32'hbf4d6bc6,
32'hbd1c1fc5,
32'h3e00cf7a,
32'h3e7ba1b2,
32'hbeab87d7,
32'hbe49c97b,
32'h3da01ccd,
32'h3fb6ddec,
32'hbf671b09,
32'hbfa1c610,
32'hbee8fd3e,
32'hbea87c02,
32'h3da5a1ef,
32'h3e47bbe0,
32'hbe50251b,
32'hbe1760e6,
32'h3d90f790,
32'h3df2eac5,
32'h3d313569,
32'hbe8a0539,
32'hbce07b1f,
32'h3d4ba556,
32'hbf66a37c,
32'hbe3ccc6c,
32'hbef71fa5,
32'h3f29aba9,
32'hbf0e4d3f,
32'hbf402bc6,
32'hbf4f42c2,
32'hbf9650fc,
32'hbf9960d9,
32'h3ed685db,
32'hbf1337b5,
32'h3ea647d4,
32'hbee5437a,
32'hbeeb1e48,
32'h3e69b4ef,
32'h3f7acf92,
32'hbeffbd18,
32'hbf9cab38,
32'h3eaa46fc,
32'hbeed774c,
32'hbddcf600,
32'hbf6614d0,
32'hbf242e5c,
32'hbf181410,
32'h3eba77b2,
32'h3f1c5760,
32'h3f6278c6,
32'h3d54997b,
32'h3d6b00c0,
32'hbd0d578b,
32'hbf71d86f,
32'hbe987c53,
32'h3d4cb245,
32'hbe9080ac,
32'h3f381b69,
32'hbe389a28,
32'hbeeb8f25,
32'hbf19090a,
32'hbf61d1e7,
32'h3f485886,
32'hbf446230,
32'hbe9f5ffc,
32'hbf30a5a1,
32'hbebd7ec6,
32'h3f1b1f0d,
32'h40080c43,
32'h3ca5fd43,
32'hbf3b5520,
32'h3eb00624,
32'hbf2626ee,
32'hbf87d89a,
32'hbfc67e55,
32'hbf57ddf1,
32'h3eed3c6c,
32'hbf027c7a,
32'hbfac1fa0,
32'hbf77af30,
32'h3eb214ee,
32'h3c87920c,
32'hbcd43348,
32'hbf79d58b,
32'hbfe35724,
32'h3e708f83,
32'h3fb13048,
32'hbedc9ff0,
32'hbd902c16,
32'hbf950e7c,
32'h3e813fab,
32'hbfee8143,
32'hbedaca80,
32'h3e301ea0,
32'hbf89d9fe,
32'hbf61ebcd,
32'hbf0a1515,
32'h3fa4d294,
32'h3f75aa3f,
32'h3f1066da,
32'hbf329afe,
32'h3ed35da6,
32'hbe6f6cb0,
32'hbe4c6ce9,
32'h3def57e7,
32'h3e1857d0,
32'h3f037cce,
32'hbe95048c,
32'hbce15033,
32'h3e136e08,
32'h3f89f9d8,
32'h3dd15ca7,
32'hbd99a64d,
32'hbdc1704f,
32'hbddf60d2,
32'hbd28bf36,
32'hbd7925f1,
32'hbd89534b,
32'hbe044fa6,
32'hbd18874b,
32'h3e599527,
32'h3a1b172e,
32'hbe446d91,
32'h3bb3ef3a,
32'hbeff1454,
32'hbeed7eea,
32'h3c3246d1,
32'hbe48500e,
32'hbe674044,
32'h3cbf9bbd,
32'h3cfb1f4a,
32'hbd49e988,
32'hbd8b387a,
32'hbd030428,
32'h3c4c7032,
32'h3cd25208,
32'h3d24d7af,
32'hbd14c1a7,
32'hbd298294,
32'h3caaa641,
32'hbd2e5c85,
32'hbd4d75f9,
32'h3d81f511,
32'hbdb7de04,
32'hbc7720e1,
32'hbc50b544,
32'h3d098303,
32'h3de4af0b,
32'h3bfddcb8,
32'h3cd91447,
32'h3dbc7f15,
32'hbe035bcb,
32'h3d326005,
32'hbd984e69,
32'hbb74ec44,
32'hbccd5299,
32'h3c5e4b68,
32'hbdba10bc,
32'h3d630de7,
32'hbd931a0f,
32'hbcc47c3e,
32'hbcd821bd,
32'h3ec95572,
32'h3e7cac3d,
32'h3e5c64d4,
32'h3e595ce9,
32'hbda870fc,
32'h3c3b8cfa,
32'h3e60148c,
32'hbeadc4f8,
32'h3ea98cc0,
32'hbd31ff54,
32'h3c141644,
32'h3f1be188,
32'hbf1ffee2,
32'hbe16cdc9,
32'hbe837e6e,
32'hbdf96650,
32'h3e74bc3e,
32'h3f821944,
32'h3f025e4f,
32'hbd5cbdbb,
32'hbe6906d2,
32'h3da99f9b,
32'hbf2ef58c,
32'hbf3b0d63,
32'h3f6dd7b4,
32'hbf185352,
32'h3ec2ea2e,
32'hbf23975f,
32'hbeefe873,
32'hbdc6a5cd,
32'h3dfdcbde,
32'hbd3283dd,
32'h3d7eb765,
32'h3d93eec3,
32'h3e8690ab,
32'h3da3cc9a,
32'h3e763c5a,
32'h3e4768de,
32'h3f1452d1,
32'hbd824fb8,
32'h3cc7f2d2,
32'h3dd2f10e,
32'hbf11e082,
32'hbf423327,
32'h3de31ed6,
32'hbdf33806,
32'hbe72fba7,
32'h3e920310,
32'hbe229ed1,
32'hbf026419,
32'hbe54aa47,
32'h3d9949e1,
32'h3e78b5dc,
32'hbf9b9abb,
32'h3ef5cedd,
32'hbe9d0860,
32'h3ed3bf17,
32'hbf024488,
32'hbec4f6dd,
32'hbbd2cf94,
32'h3f45732f,
32'h3ec7a605,
32'hbf422f59,
32'hbe4b40fa,
32'h3f01f3a2,
32'hbf84a801,
32'hbd1812e6,
32'h3e347e4a,
32'hbf142e52,
32'h3d1c1b6d,
32'h3cc40d59,
32'hbfb1bfcf,
32'hbf71812f,
32'hbf2e1838,
32'h3da0e310,
32'h3e099010,
32'h3e38621d,
32'h3edb346e,
32'h3ea55087,
32'hbf3ce91c,
32'hbeddeadb,
32'hbe7a1395,
32'h3c8ff1d7,
32'hbe202389,
32'h3e47d5e2,
32'hbeef4b36,
32'h3e1b0e63,
32'hbdf6087a,
32'h3f0668b1,
32'h3e807113,
32'hbd42f6cf,
32'h3f19d820,
32'hbe181845,
32'hbf028b9b,
32'h3dd873f9,
32'hbf372a93,
32'h3d222b14,
32'hbec8c9a7,
32'hbe2037ee,
32'hbd8d6664,
32'hbd538dc5,
32'hbf2d5e27,
32'hbfd69123,
32'hbf0bdcb4,
32'h3e2945a1,
32'h3f5804bf,
32'hbebc27d1,
32'h3e832c6a,
32'hbee40bef,
32'hbf717654,
32'h3e935729,
32'hbe9b12d4,
32'h3e944169,
32'h3cef2631,
32'hbea6060d,
32'h3ea70609,
32'hbf97b722,
32'hbf717988,
32'hbef9f5d8,
32'hbf14bbce,
32'h3e09e573,
32'h3ed1c041,
32'hbeeaf531,
32'h3c7f1565,
32'h3e7476e2,
32'hbe810a9f,
32'h3dbac7ee,
32'h3f008c01,
32'h3ed8d9ee,
32'hbdd967a4,
32'h3cf145ba,
32'hbecc01dd,
32'hbff65695,
32'hbf3f7241,
32'h3e000a31,
32'h3f364d94,
32'h3e778fb3,
32'h3e81a6c9,
32'hbcac3aec,
32'hbf629428,
32'hbde682a2,
32'hbf05bb52,
32'hbd8c9cad,
32'h3e562e4e,
32'h3eac6275,
32'h3d3e4a5f,
32'hbf2284d2,
32'hbfc6e1e6,
32'h3e3b1b0e,
32'hbe220b38,
32'h3e280115,
32'h3e25139f,
32'h3ea8a936,
32'hbdf9b501,
32'hbe33a1f2,
32'hbf619e49,
32'hbe5ab8c9,
32'hbdff0f9e,
32'hbe86b98b,
32'hbd3f57cc,
32'hbd89827c,
32'hbea7d16e,
32'hc00ac34b,
32'hbf1df54d,
32'hbdaf71df,
32'hbef0bdd2,
32'h3e4582aa,
32'h3e08205a,
32'hbe597a3d,
32'hbe0d774a,
32'hbcc68c68,
32'hbd83018c,
32'h3d8f3930,
32'hbfb4e075,
32'hbf0cd52c,
32'hbd14e893,
32'h3d9a7b0d,
32'hbfc31de5,
32'h3d401f94,
32'hbf72d036,
32'h3e39df1f,
32'h3d364043,
32'hbd08d5c6,
32'hbde63c44,
32'h3eb28abd,
32'hbf645144,
32'h3ed6c289,
32'hbe0d9b4b,
32'h3d0bb4e9,
32'h3d17270b,
32'h3c6f75df,
32'hbe66bdc0,
32'hc007445e,
32'hbf7b3e13,
32'h3d9c8c11,
32'hbf5442b5,
32'h3b1a3c86,
32'h3d268578,
32'hbdcfeecf,
32'h3d4f7b6e,
32'h3d2c0b0c,
32'hbf0bb725,
32'hbe3362ec,
32'hc00564ca,
32'h3e261aa9,
32'hbdbe2abb,
32'hbdb629a4,
32'hbf131065,
32'h3d376519,
32'hbf8919e1,
32'h3dbd2221,
32'h3f0b15bf,
32'hbecb2b2a,
32'hbd85027b,
32'hbe2aed44,
32'h3dc4e638,
32'h3ef1f3d9,
32'h3d33efa1,
32'h3d5c413e,
32'hbcefb4a4,
32'h3c35ddbc,
32'hbd6bc1b0,
32'hc000d59c,
32'hbcaba31c,
32'h3e04d861,
32'hbf8abccc,
32'hbe08eac9,
32'hbddc975f,
32'h3e80c6d0,
32'h3e238231,
32'h3e1a3eb9,
32'hbc42d944,
32'h3d7bfe55,
32'hc0608a6f,
32'hbd6de9ed,
32'hbe164fb5,
32'h3dfd7aad,
32'hbef8a761,
32'h3ee5420e,
32'h3d8496b0,
32'h3dad3d59,
32'h3dca4db3,
32'hbd8e9059,
32'hbdb304d2,
32'hbd654666,
32'h3f002917,
32'h3e3b934c,
32'hbdbc5940,
32'h3dd9d415,
32'h3d21fdd6,
32'hbdf1c207,
32'hbe29950e,
32'hc006d973,
32'hbe17cddf,
32'hbddfc2b9,
32'h3d1249f3,
32'hbd2cd684,
32'hbdde037b,
32'h3e89b3fd,
32'h3d2aeaf3,
32'h3e5ee10f,
32'hbe2ea458,
32'h3e293e01,
32'hc044f63e,
32'hbece4e28,
32'hbcd11e96,
32'h3d88f9e1,
32'hbe69fc0b,
32'h3e4bc48a,
32'hbe15b6ed,
32'h3ddf54fe,
32'h3d2a2bbc,
32'h3d8273cb,
32'h3d6d71f4,
32'h3e07388b,
32'h3f2b4ff7,
32'hbcf2f5c6,
32'hbf1f4849,
32'h3d9cc8ec,
32'hbcc4ebd2,
32'hbdd17e31,
32'h3e3d6a1c,
32'hbf73fbdc,
32'hbd3ddc64,
32'hbe425d15,
32'hbe3836fe,
32'h3dfb55e2,
32'hbd7b627f,
32'hbdc95431,
32'h3e791eda,
32'h3e10f2a5,
32'hbe602aa7,
32'h3c08ac59,
32'hbf8f8e0c,
32'hbe098418,
32'h3db00bb4,
32'h3e3245f0,
32'hbe9210ab,
32'h3decea6d,
32'hbf32d579,
32'h3e8e4033,
32'hbf41930d,
32'h3e954815,
32'hbe0fe022,
32'h3e2fc8f5,
32'h3e75fb11,
32'h39eee38a,
32'hbed15a3e,
32'hbeba72b5,
32'hbc431811,
32'h3d65391f,
32'hba0fa85b,
32'hbf8ee522,
32'hbee1b1bc,
32'hbe3c70e7,
32'h3a1baf11,
32'h3ec403b2,
32'h3e3b05b9,
32'h3dc0ee7c,
32'h3e896f76,
32'hbd66fc99,
32'h3d41f937,
32'h3e27c2ed,
32'h3b80ce14,
32'h3e1ff73b,
32'h3d99fae8,
32'h3d785394,
32'hbd2b4546,
32'h3e56be2a,
32'hbd4906c7,
32'h3e0faecc,
32'hc0220d34,
32'hbd0a8f80,
32'hbe658f0e,
32'h3e822208,
32'h3e8c1e7b,
32'h3e0ed90f,
32'hbdfbc9b0,
32'h3d01ebb0,
32'hbc351759,
32'h3bac5470,
32'hbe86d196,
32'hbf33c752,
32'hbf433447,
32'h3c6299a1,
32'hbf063352,
32'h3ec94a97,
32'hbdf0700a,
32'h3d7eb2eb,
32'h3ed4622f,
32'hbd8dd149,
32'hbd3d7b26,
32'hbc572dd8,
32'h3e5b6b98,
32'hbed7a89f,
32'h3d87aabc,
32'hbe24e891,
32'h3e2d7443,
32'h3ebe3a32,
32'h3d88c0fa,
32'hbf230d78,
32'hbf9fa641,
32'hbe982d57,
32'hbe2bea8c,
32'h3ea399a6,
32'hbd01b172,
32'h3e87fa83,
32'hbea4226b,
32'h3e589534,
32'hbe06bac9,
32'h3ca5b9a1,
32'h3c3d90ba,
32'hbf10cedb,
32'hbf6f1cad,
32'h3cc3c5d0,
32'hbee8d9f9,
32'hbf0b708c,
32'hbf2c3323,
32'hbdb9b50e,
32'h3eac1c7b,
32'hbde50b8d,
32'h3e1bbe8a,
32'hbe081275,
32'h3e956540,
32'hbfc6abc0,
32'h3e089df8,
32'hbe172004,
32'h3ded886b,
32'h3e00a732,
32'h3e9fc3a9,
32'hbeba68bb,
32'hbeb826f7,
32'hbf5d5a6e,
32'hbec2f747,
32'h3e7b1e91,
32'h3e374dd5,
32'h3e972b23,
32'hbd0eaf4f,
32'h3d4a523a,
32'hbdd6cb9d,
32'h3c96608d,
32'hbd9f1892,
32'hbe84f62c,
32'hbf4264a9,
32'h3e55da35,
32'hbe976281,
32'hbef7c456,
32'hbe3348c1,
32'hbf3558ab,
32'h3d82e1e7,
32'h3b841a68,
32'hbdf0042f,
32'hbe9b463f,
32'h3ea63f7d,
32'hbe57c9f5,
32'h3db46262,
32'hbf20d1cd,
32'h3d9a1583,
32'hbe81ace7,
32'h3e573d9c,
32'hbf414ba3,
32'hbe9ea18c,
32'hbf8c5890,
32'h3a8a38e1,
32'h3e80ff26,
32'hbd541201,
32'h3e91a24e,
32'hbe80e2d3,
32'hbb719b53,
32'hbd103c39,
32'hbd25bf1b,
32'hbeea9fe2,
32'hbf4c24a2,
32'hbf135ec5,
32'h3e898c2b,
32'hbd835944,
32'h3cebed3d,
32'h3f0e2582,
32'hbf42c87b,
32'h3e588fe6,
32'h3ec44061,
32'hbe2f5f1d,
32'hbe4cf2fb,
32'h3e52d86d,
32'h3e432fb1,
32'h3cbbef96,
32'hbf22a8e7,
32'hbe9a3a7f,
32'hbe1a8497,
32'h3e8ab95b,
32'h3e18c14b,
32'hbca49229,
32'hbf655b6b,
32'h3e08fd50,
32'h3dc17893,
32'hbe945d3b,
32'h3e69075c,
32'hbdc717a1,
32'h3e186d3d,
32'hbdca2561,
32'hbc900331,
32'hbe7ce80e,
32'hbdfeb872,
32'hbebac392,
32'h3d1508f3,
32'h3e8965bc,
32'h3dae97c3,
32'h3e79e753,
32'hbe9cc041,
32'h3e302dca,
32'hbda6079a,
32'hbea5b0d6,
32'hbe32db2b,
32'h3eae6cc6,
32'h3df4317e,
32'h3d8b2539,
32'hbfc65c19,
32'h3d91d26b,
32'hbdcac83d,
32'h3dee7d07,
32'hbcdc6ce5,
32'hbd1699d7,
32'hbf3eb775,
32'h3e58bf4b,
32'hbe2f50c8,
32'hbe0d07ca,
32'h3ea2726b,
32'h3c3f69b4,
32'hbe3febc7,
32'hbdb1189e,
32'h3d8bdd31,
32'h3e945935,
32'hbe7bf373,
32'hbec6055e,
32'h3e228f0c,
32'h3e07795d,
32'hbda4ff62,
32'h3e733ae7,
32'h3e496868,
32'h3d3d3edc,
32'h3dbb064f,
32'h3e931c22,
32'hbd37261b,
32'hbc6fc9f1,
32'hbede5f4e,
32'h3cb877db,
32'hbfd15935,
32'hbea05241,
32'h3e079b40,
32'hbe6918ae,
32'h3e1a9f9b,
32'hbe52c5a3,
32'h3d702df9,
32'h3e37ca31,
32'hbd2ae6e3,
32'hbe1af724,
32'h3eb0105d,
32'h3e72c348,
32'hbed92619,
32'hbd0eb2ea,
32'h3d84e6fc,
32'hbe2cc102,
32'hbe9c676d,
32'hbeab5a1f,
32'h3db0cbd3,
32'h3e2fce8c,
32'h3e0defb4,
32'h3e6d9619,
32'h3e242db8,
32'hbdc94a13,
32'h3e4a4bfd,
32'h3deedbdd,
32'hbe9aef47,
32'h3e145421,
32'hbe36771a,
32'hbd5911a8,
32'hc003043f,
32'hbdcde248,
32'h3d0bd899,
32'hbe9866df,
32'hbe5ce811,
32'h39761eb5,
32'h3e40b52c,
32'h3de70957,
32'hbf38d45b,
32'hbf14ef09,
32'hbd971035,
32'hbe3d778d,
32'hbf848c5e,
32'hbe2fbaa9,
32'hbd6fdc17,
32'h3df90c7e,
32'hbd184999,
32'hbefb0836,
32'h3e4c89b5,
32'h3dace2e9,
32'hbd0bb47b,
32'h3c51b12a,
32'h3d883002,
32'hbdc6e536,
32'hbdc1618a,
32'hbf09f18a,
32'hbe16b3b0,
32'hbe589f79,
32'hbde3686e,
32'hbdee7c5d,
32'hc015a583,
32'hbea3be14,
32'hbef08f12,
32'hbf10f496,
32'h3dea6d0b,
32'hbe089d17,
32'hbe0d727d,
32'hbdf2351b,
32'hbf44c6ba,
32'hbdc02ee5,
32'h3e4657fb,
32'h3dff9dbf,
32'h3e14ec99,
32'hbe01e065,
32'hbc15924b,
32'hbc80793c,
32'h3dc836f2,
32'h3ce45c81,
32'h3e049763,
32'hbee513e0,
32'hbea2e397,
32'hbd9a94ce,
32'h3c398e3e,
32'h3cbcc3dc,
32'hbc318712,
32'hbe96eaef,
32'h3d81e02d,
32'hbdcbe2da,
32'hbe44dde8,
32'hbca73f95,
32'hbfbc785a,
32'hbe9783c4,
32'hbeb9eb37,
32'h3ec645cf,
32'h3e1e8d0c,
32'h3bc4b0ad,
32'h3e75fbed,
32'h3cbb6e53,
32'hbfa2dafc,
32'hbe54066c,
32'h3e988695,
32'h3e2a895f,
32'hbd9eab1e,
32'hbe0e8a14,
32'h3d5c0276,
32'h3e087e9f,
32'h3e062fa2,
32'hbda24511,
32'h3d542ced,
32'hbf2031e3,
32'h3dbf5089,
32'h3db7e2e6,
32'hbd05972f,
32'h3c0e4bd8,
32'hbe451535,
32'hbeabf785,
32'h3c42beae,
32'hbe9f56fa,
32'hbec06ca4,
32'hbdb854e4,
32'hbf69bf55,
32'hbe1dacef,
32'hbefbb984,
32'h3dc6112f,
32'hbe0f4ae3,
32'hbb6325a6,
32'h3e54fdfc,
32'h3e94a10e,
32'hbf7a7582,
32'hbf628da4,
32'hbde3f273,
32'h3d787f0f,
32'h3ea2480b,
32'hbd269a98,
32'hbd60a08b,
32'h3c68ab2d,
32'h3db6a737,
32'h3db35278,
32'h3edb276a,
32'hbfb2e6fb,
32'h3ea85be1,
32'h3e9b02ae,
32'hbd3ff45c,
32'hbd80fbc7,
32'hbd88ab44,
32'hbf13b0b4,
32'h3e92dcbb,
32'hbf161f5d,
32'hbe62ef57,
32'hbf024bcf,
32'hbf20a31c,
32'hbe8682e1,
32'hbf2331bc,
32'hbf201ced,
32'hbdcbd605,
32'hbef8cde9,
32'h3f015874,
32'hbd02b3d8,
32'hbf2cd452,
32'hbe8071fb,
32'hbeb516ad,
32'hbea70f6a,
32'h3ee0c839,
32'hbc93264f,
32'h3ca3acef,
32'hbd4343db,
32'hbe563ad8,
32'hbea5ec73,
32'h3f3bdcca,
32'hbf40afb5,
32'hbe4c8151,
32'h3edc5b14,
32'hbf065d80,
32'h3e017c48,
32'hbe199019,
32'hbe523942,
32'h3ee3c8b3,
32'hbdd45efe,
32'hbf7e1d85,
32'hbe8dc992,
32'hbf2168b5,
32'hbe9aab6f,
32'hbecf911e,
32'hbedc0987,
32'hbe9e8610,
32'hbce685db,
32'h3eb815be,
32'hbfaa7892,
32'h3ae98daf,
32'h3f5c5cb3,
32'hbea88313,
32'h3ef390d5,
32'hbe70e708,
32'h3c40d889,
32'hbbcfaab6,
32'h3e11e0b5,
32'h3e64bf39,
32'hbe58f7e2,
32'h3f102dfd,
32'hbf37c50d,
32'hbda434c0,
32'hbf6cb5d0,
32'hbf1450e6,
32'h3da7faec,
32'h3e577382,
32'hbf1de895,
32'h3eb12e4e,
32'hbb3ba696,
32'hbf8d91dd,
32'hbee10af7,
32'h3f3de3b3,
32'h3c73e57d,
32'hbe5ae247,
32'hbe6ec10d,
32'hbf1c270a,
32'h3d881f9e,
32'hbeb90a7e,
32'hbe2f47d8,
32'hbee6806c,
32'h3f9fc16a,
32'h3e93c76a,
32'h3f7929a7,
32'h3e415953,
32'hbd2f360b,
32'hbcaaf870,
32'hbed78e98,
32'h3e501f4f,
32'h3f062c60,
32'h3e0247e8,
32'hbedd8b54,
32'h3f5bd6db,
32'hbe88ee6d,
32'h3f47735e,
32'h3f18cab9,
32'h3f0839e1,
32'hbf5166f1,
32'h3d9b1ea4,
32'h3f89b2e3,
32'hbd26b9cb,
32'h3ed9afcf,
32'h3f770201,
32'h3fc17f7d,
32'h3dc211de,
32'hbf971c8c,
32'hbea965bf,
32'h3ef8ddd6,
32'hbf326388,
32'h3eb678d8,
32'hbe03bc01,
32'hbf15680b,
32'h3e98d514,
32'hbcebae5a,
32'hbdeec956,
32'h3cd90f6c,
32'hbcd84e45,
32'hbfc7ebbc,
32'h3edaae6a,
32'h3fa8890a,
32'h3f37bef1,
32'hbed2e530,
32'hbe294190,
32'hbf480134,
32'h3f0543b6,
32'h3bbfd0b1,
32'h3f28ee35,
32'hbf9ead19,
32'hbf49d217,
32'h3e72a948,
32'hbc7abd23,
32'h3ed0aa46,
32'h3f0a15b6,
32'h3fc73118,
32'hbde1dcf5,
32'h3c8b5a16,
32'hbda41b9e,
32'h3d8885c7,
32'h3daae1bb,
32'h3d470d55,
32'h3f1777f5,
32'hbe8c6c13,
32'h3e7c64cd,
32'h3f6caab5,
32'h3f8afc56,
32'h3d209637,
32'hbc771f16,
32'h3dc43496,
32'hbe1301e5,
32'h3d008331,
32'h3db0bc23,
32'hbdcc8c0a,
32'hbeb2cc9e,
32'hbcc3d9d9,
32'h3d0c1dd8,
32'hbe45563a,
32'hbef36c70,
32'hbde2d3d0,
32'hbf5c668f,
32'hbf07ba11,
32'h3d36dd8c,
32'hbe780550,
32'h3d3dd175,
32'h3f05b221,
32'hbe879e95,
32'hbdd0b1f5,
32'hbc920122,
32'hbd2893a5,
32'h3c5c5655,
32'hbcb22530,
32'h3d103cbf,
32'h3d1379bd,
32'hbcffce25,
32'h3d2ee900,
32'hbe0236bf,
32'h3d5785e1,
32'h3d9c0c9a,
32'h3ba11639,
32'h3da30ebb,
32'hbde727e2,
32'h3da5f9fa,
32'h3c0a1106,
32'hbddf1a0e,
32'h3ca44bc9,
32'hbdd50055,
32'hbc0a44aa,
32'hbd65f3c9,
32'hbc2b88f8,
32'hbd32bd93,
32'h3cb0084e,
32'h3b28bbe3,
32'h3cc21598,
32'hbdbf6262,
32'h3c3e8d70,
32'h3d123372,
32'hbbda863e,
32'hbd6d9089,
32'hbddd5c77,
32'h3e3e44cb,
32'hbd6fe74c,
32'hbd151fdb,
32'hbde4e3cc,
32'h3e7949e5,
32'hbd6ff9ed,
32'h3d08adc3,
32'hbccb8456,
32'hbdb694aa,
32'h3f112bad,
32'hbf084fae,
32'hbd879031,
32'hbe6b7e4e,
32'hbdeb4061,
32'h3f014950,
32'h3f17bd67,
32'h3e944c19,
32'h3d34947e,
32'hbe321d87,
32'hbd948e78,
32'hbdff8c09,
32'hbf0cfbf1,
32'h3e009a67,
32'hbe58d155,
32'h3da05ad5,
32'hbf0eb74a,
32'hbe51451e,
32'hbea7e60b,
32'h3f2ed213,
32'h3e5075d8,
32'h3e434833,
32'h3cda67e0,
32'hbe6d1787,
32'hbf1760cd,
32'h3d4254fa,
32'h3ee86626,
32'h3d65dca5,
32'hbda051ff,
32'hbd12986e,
32'hbf5bd4a7,
32'hbeb54753,
32'h3e864fa2,
32'hbc59ec03,
32'h3eb2494b,
32'hbe79da5c,
32'h3eda6c1f,
32'hbe2b8c78,
32'hbf647884,
32'h3ebfb61e,
32'hbdeff15f,
32'hbf15facb,
32'hbee5945c,
32'h3f72e8d4,
32'h3e2e850a,
32'h3e8dfe70,
32'hbf0c4cee,
32'hbf8679f4,
32'h3e32c15d,
32'hbdd237f7,
32'h3f62ffef,
32'hbf01230a,
32'hbd6f9c6c,
32'hbe2899aa,
32'hbcf1d1dc,
32'h3fadd265,
32'hbf0b11f6,
32'hbe398f30,
32'hbd008421,
32'h3d5a3906,
32'hbfad08aa,
32'hbf484d24,
32'hbf511c31,
32'hbdc2dd64,
32'h3f297a92,
32'h3cfb33b4,
32'hbd91c2fe,
32'hbf0d146d,
32'hbf43126f,
32'hbe1921ea,
32'hbf04ad29,
32'h3dd49505,
32'hbf80142d,
32'h3c737cff,
32'hbedf0bc7,
32'h3d8ff07e,
32'hbe11240c,
32'h3f134ff7,
32'h3e158449,
32'hbee817b9,
32'hbe4a4458,
32'hbcccff0e,
32'hbe6347c6,
32'h3e351786,
32'h3e9529ba,
32'h3f197817,
32'hbe98e94b,
32'h3ebf604f,
32'hbdbe50e0,
32'hbd3ec202,
32'hbe8fa5bc,
32'hbfa5b051,
32'hbf80dbd0,
32'hbd32256a,
32'h3e1820b7,
32'h3d2dcea7,
32'h3ed054f1,
32'hbe846141,
32'hbf97001d,
32'h3e236d5d,
32'hbefca43d,
32'h3f0376e9,
32'hc007257b,
32'hbea4fe6b,
32'hbf1185b0,
32'hbf943bd3,
32'hbf08b304,
32'hbdc4eab2,
32'hbfadffbb,
32'hbd3e4ca1,
32'h3e969c7b,
32'hbdcb52d5,
32'hbebbd1c3,
32'h3dc59881,
32'hbd913194,
32'h3ef0d629,
32'h3ee54d19,
32'hbeb53461,
32'hbd17b60e,
32'hbda35fcb,
32'hbe1c7ca7,
32'hbf9876b4,
32'hbf28a357,
32'hbe0108a4,
32'hbebb7450,
32'h3d98b481,
32'h3e0b84fd,
32'hbcf38028,
32'hbf192dc7,
32'h3d90a02f,
32'hbef1bdc9,
32'h3e49df24,
32'hc0117547,
32'h3d83e78c,
32'h3dbf5fb4,
32'h3e293722,
32'hbeaa2c54,
32'h3e657d8c,
32'hbfcf7783,
32'h3c24d581,
32'h3e29a166,
32'h3ec33e3a,
32'hbda19759,
32'hbd4a12d9,
32'h3e754880,
32'h3d105824,
32'hbee49915,
32'h3eaf17dd,
32'hbd24a63c,
32'hbd83a092,
32'h3dbc2802,
32'hbf7bee42,
32'hbfb197cc,
32'hbef82a10,
32'hbf9556d1,
32'hbdba362c,
32'h3db42dfc,
32'hbcb146af,
32'h3e695110,
32'hbd115d02,
32'hbe7f00ce,
32'h3c299ba2,
32'hc0189545,
32'hbd58e855,
32'hbe75edcf,
32'h3ecd5f08,
32'h3f0e65a8,
32'h3e88fee5,
32'hbeed151f,
32'h3d760719,
32'h3d356c20,
32'h3e876d43,
32'h3df391ef,
32'h3e6580ea,
32'h3ea97f8c,
32'hbea9f788,
32'hbf33efec,
32'h3f0ce86f,
32'hbdc4f5af,
32'h3cb50e6b,
32'h3e59ba8f,
32'hbf3e9751,
32'hbfb40cba,
32'hbe570d68,
32'hbf51114c,
32'hbda4be59,
32'h3e3b3d65,
32'h3ca7ff81,
32'hbd363b10,
32'h3d5120d0,
32'hbe7b83ea,
32'hbbf8aa2f,
32'hc03546a1,
32'h3ecbf06f,
32'hbdbcabbc,
32'h3de9369a,
32'h3efed9bf,
32'hbec1e006,
32'hbe9fb689,
32'h3e07e22e,
32'h3dcad83b,
32'h3ddd0e4e,
32'hbe0e8ded,
32'h3d0e3a61,
32'h3edb5984,
32'h3c484078,
32'hbf8c3d39,
32'h3cd7caa7,
32'hbd159780,
32'h3cb25165,
32'h3e22eb1f,
32'hbe7769d5,
32'hbfb4955b,
32'hbe835450,
32'hbf903496,
32'h3e27289e,
32'h3deb4432,
32'h3e518028,
32'hbd749f14,
32'hbdaca646,
32'hbd44f92b,
32'h3e3b9b3e,
32'hbf822d69,
32'h3f35f1ed,
32'hbd898cd2,
32'h3e49c489,
32'h3e1f2cc4,
32'h3ed49733,
32'hbf4f571a,
32'hbda19071,
32'h3e315b2c,
32'h3e2336c1,
32'h3d6288b7,
32'h3c9a8aa4,
32'h3eef3278,
32'h3dc62fff,
32'hbf46a84c,
32'h3e25f07f,
32'h3c1f4a53,
32'hbcbd6715,
32'hbde1b062,
32'h3d3744d4,
32'hbf994d23,
32'hbed606d1,
32'hbf2f448d,
32'h3de51a84,
32'h3c88f984,
32'hba2a2fd3,
32'h3e126e5e,
32'hbe38a20b,
32'hbdd9e3fb,
32'hbdecca67,
32'hbc59c927,
32'h3db6be3b,
32'h3e3db8ce,
32'h3c620ee7,
32'h3ecc76c4,
32'h3c92f03c,
32'hbf37fb75,
32'h3e47c5c1,
32'hbf7be0ad,
32'h3ef222d3,
32'hbe8291bd,
32'h3e06be8b,
32'h3c8440fd,
32'hbd968fe4,
32'hbf546223,
32'hbe507a07,
32'hbd92de9a,
32'h3d05f905,
32'h3d5c8db7,
32'hbe694c7f,
32'hbfd37a18,
32'hbe83117e,
32'hbe6bc85d,
32'h3ee30d03,
32'h3b69db52,
32'hbd1b2c81,
32'h3eec691a,
32'hbc05aa08,
32'hbd08e478,
32'hbe2ae26c,
32'h3e2874e5,
32'h3ed911bd,
32'hbe1513e2,
32'h3e94a06d,
32'h3e274590,
32'h3ebef24d,
32'hbdfb8c62,
32'h3da0ba4f,
32'hc033b9c2,
32'h3d3b4534,
32'h3d8d2c34,
32'h3e8459ac,
32'hbe1897ab,
32'hbe70555b,
32'hbeb00902,
32'hbec1d430,
32'hbcc8133c,
32'hbcf9f5fe,
32'h3d5d4dc1,
32'hbdbbea63,
32'hc0102689,
32'h3e2001d7,
32'hbf0bf907,
32'h3eb734a7,
32'h3de01d33,
32'h3e678f58,
32'h3e91d40c,
32'h3e4b5b39,
32'hbe2c1125,
32'hbda53094,
32'h3e312269,
32'h3ef8dae8,
32'h3e8e0716,
32'h3e7a10c7,
32'h3eaa7d96,
32'h3ec10705,
32'hbece0194,
32'hbeb1fa64,
32'hbf477336,
32'hbeedaa18,
32'hbeabb273,
32'h3ea00b78,
32'hbe25d28f,
32'h3d3e25ce,
32'hbea168af,
32'hbe286dcc,
32'h3c78c696,
32'h3c9a1525,
32'h3bd2cf09,
32'h3e0ad1e7,
32'hbfe84bd0,
32'h3e802304,
32'hbe888c40,
32'hbd930f7a,
32'hbe934af4,
32'h3de90d5b,
32'h3ec81a04,
32'h3e070efd,
32'h3e433e0d,
32'hbe80db55,
32'h3ebd7c4e,
32'hbf357bbd,
32'h3db9f064,
32'h3e40f7c9,
32'h3eb11393,
32'h3c250201,
32'h3e7db574,
32'hbf76180b,
32'h3ea3e496,
32'hbf73e037,
32'hbef2b3ba,
32'h3df9ad44,
32'h3e2224df,
32'hbdbcba6d,
32'hbe0ce9e4,
32'hbeae9df5,
32'hbcc0d738,
32'h3d07a61b,
32'h3a76f7ca,
32'h3cecf3ed,
32'hbfa2dc0e,
32'h3d892103,
32'h3c5dea5f,
32'hbefc71a2,
32'hbe4f57c6,
32'hbe0d4968,
32'h3e033019,
32'h3e0b036d,
32'h3e2bc8a7,
32'hbe5024d6,
32'h3ee0bbcd,
32'hc001546f,
32'hbccf2146,
32'hbd262641,
32'h3ecb2d1f,
32'hbe6a8e0a,
32'h3e2fccae,
32'hbf3654e8,
32'hbe9235dd,
32'hbfb6b8a3,
32'h3cbff4c1,
32'h3db0526d,
32'h3ea63ecd,
32'h3e37dc2a,
32'hbd6a2711,
32'h3dc9bb71,
32'hbd8864dd,
32'h3cd20e3d,
32'hbe3f4cd9,
32'hbf1150f6,
32'hbf76b89c,
32'h3e6d971f,
32'hbe06360d,
32'hbe999718,
32'hbd4b2879,
32'hbec5991b,
32'hbcc6cf72,
32'h3d6fa05a,
32'hbe18e979,
32'hbe2dba2c,
32'h3d5ff8a6,
32'hbea06c9d,
32'h3da87aa5,
32'h3d1a03e9,
32'h3e3645dc,
32'hbee7f62e,
32'h3e281a1b,
32'hbf1e12c0,
32'hbe00fdaa,
32'hbfa8a4dd,
32'hbc95bd09,
32'h3d886b8b,
32'hbd7c1005,
32'h3e50ddf9,
32'hbbc1a619,
32'hbdb61734,
32'h3cb150a5,
32'hbcfb7ecc,
32'hbe0830c6,
32'hbf013b4e,
32'hbec0dc67,
32'h3e806d7e,
32'hbdd49561,
32'hbd62c459,
32'h3e9c473e,
32'hbf451ae1,
32'h3e29723f,
32'h3cdfc017,
32'hbd8471df,
32'hbe26eba0,
32'hbe28e7a8,
32'h3dad1b6a,
32'hbe016e7f,
32'hbeacc97a,
32'hbdba8f8c,
32'hbe308894,
32'h3dc33895,
32'hbdb19f62,
32'hbe1919d4,
32'hbfa7879e,
32'h3e102b93,
32'hbe61f4df,
32'h3d567fce,
32'h3e807784,
32'hbec69257,
32'hbd16ac1b,
32'hbdf5d0cd,
32'h3c3e99f7,
32'hbc64e9b7,
32'hbe2c56c9,
32'hbedf5d37,
32'h3da7a2f8,
32'h3d3df293,
32'hbcb153e6,
32'h3eb3e980,
32'hbe504424,
32'h3e99175b,
32'h3d072943,
32'h3d430ba2,
32'hbd769f0f,
32'h3e113358,
32'h3deafea5,
32'hbdec47cc,
32'hbefcd3ab,
32'h3e15c60e,
32'hbd729589,
32'h3d36b2e4,
32'h3da830ec,
32'h3d131c7f,
32'hbea9f957,
32'hbcca7716,
32'hbd4fc3dc,
32'hbc1a4689,
32'hbd5530f1,
32'hbd3590d8,
32'hbec98fd3,
32'hbd79c08d,
32'h3d0a9e7f,
32'hbc6fcd55,
32'hbea80c45,
32'hbeb5d95b,
32'h3ddbb96c,
32'h3e78479a,
32'h3d8f05ad,
32'h3ed9e5be,
32'h3ebaf9ee,
32'h3da17d25,
32'h3cb5c8d2,
32'h3e34c025,
32'hbe44e26f,
32'h3e2459c3,
32'hbe6cdacc,
32'hbe3cf11c,
32'hbf2bee22,
32'hbe08b360,
32'h3e94abd6,
32'hbedbda74,
32'hbdae01ba,
32'hbd4d7c38,
32'hbe1ee525,
32'hbe4e8166,
32'hbd8d6172,
32'hbe2e1440,
32'hbce72fab,
32'hbd84c2db,
32'hbf7552d1,
32'hbe0cd8dd,
32'hbd0c4aa0,
32'hbcf6fe21,
32'hbc758bed,
32'hbec05ebd,
32'h3de2c3ec,
32'h3e90af76,
32'h3d9b3f71,
32'h3e4a0fad,
32'h3e268a3d,
32'h3caab0d7,
32'h3e14c2a8,
32'h3e4d87b1,
32'h3dcf7723,
32'h3d6685c6,
32'hbe7839f9,
32'hbced93fe,
32'hbfa6a579,
32'hbd7871ae,
32'hbdb46764,
32'hbe880128,
32'hbecb62ad,
32'hbe2de7f6,
32'hbe7318e1,
32'h3e4b0a57,
32'hbee5e627,
32'hbf070c75,
32'hbdb84737,
32'h3c68d2e8,
32'hbd141ec7,
32'h3c720b45,
32'hbd8ab896,
32'h3e0aefef,
32'h3da417e2,
32'hbcb41fbe,
32'h3d48d3ec,
32'h3e28e844,
32'h3d0f117d,
32'hbe2499b2,
32'hbe0da05c,
32'h3d5bd6d2,
32'h3df0cc6f,
32'h3e130dbf,
32'hbdb8e1ba,
32'hbf0fb7d8,
32'hbf2367b8,
32'hbbe5b438,
32'hbfdc396e,
32'hbe9ac5c4,
32'hbe47ffc7,
32'hbeb739aa,
32'hbd7ac2b6,
32'hbe73a96d,
32'hbe899258,
32'h3e470449,
32'hbe4a5ee8,
32'hbe3d27b1,
32'hbe183f58,
32'h3d2516a2,
32'h3e6140ff,
32'h3c04001f,
32'h3d50e6d4,
32'h3c01022d,
32'hbe68a061,
32'hbe7f95c8,
32'h3dc48f73,
32'hbf84462a,
32'h3d99fcf3,
32'hbc95d39e,
32'hbe44351a,
32'h3f26e969,
32'h3e57d942,
32'hbcc9d777,
32'hbd588ac5,
32'hbebe544e,
32'hbebf2c2c,
32'h3dc5ad36,
32'hc006b338,
32'hbe5f6a02,
32'hbe3dac82,
32'h3f24881e,
32'h3e5028f7,
32'hbd18ae3c,
32'h3dd2f49a,
32'h3d1d5a15,
32'hbe4b745f,
32'hbe05ee5f,
32'hbe47bd73,
32'hbf12a7cb,
32'hbe6d2a79,
32'h3d28dc61,
32'hbc56b029,
32'h3e967a40,
32'hbe62ea11,
32'hbdc9354b,
32'h3e061450,
32'hbfb46d2b,
32'h3ef7b3a0,
32'h3ebdde8e,
32'h3d64f703,
32'h3dd1d21c,
32'h3e9c659d,
32'h3e770d12,
32'hbda489a2,
32'h3eb7fdac,
32'h3d7bdb71,
32'h3d8726e7,
32'hc037a402,
32'h3d847c00,
32'hbe7dd029,
32'h3e645e67,
32'hbeca1aa2,
32'hbecc0240,
32'h3e05a5b1,
32'h3e6b478a,
32'hbf00149c,
32'hbeee90c4,
32'hbeb8db2f,
32'hbf00941d,
32'hbf3ddea1,
32'hbd7df89c,
32'hbd08aa9d,
32'h3e66dbdf,
32'hbcc66a54,
32'h3d1cf724,
32'h3e515960,
32'hbfab1d62,
32'h3d5b305a,
32'h3c1571d0,
32'hbecc6472,
32'hbe453921,
32'h3ea05075,
32'h3d80c320,
32'h3f1ffb9f,
32'hbcaa4ada,
32'hbf183943,
32'hbf0e41a0,
32'hc01b3c81,
32'hbcf6be1e,
32'hbd55d867,
32'h3e39af21,
32'hbf11fcd6,
32'hbe79775b,
32'h3eeb7f7d,
32'hbe71540b,
32'hbf13bac5,
32'hbe52fd8b,
32'hbf23952a,
32'h3dabb963,
32'hbf834d3c,
32'hbb413dd6,
32'hbdc0b377,
32'h3f1f3016,
32'hbe090400,
32'hbe06b9ab,
32'h3ecfc59b,
32'hbf47f1f0,
32'hbe2ff95a,
32'hbf3067f6,
32'hbf5fdbc6,
32'hbb39c38b,
32'h3d778672,
32'hbf408360,
32'h3f357be4,
32'h3e5c3d8f,
32'hbf2a431c,
32'hbeda3ee6,
32'hc004cfe6,
32'h3ee66e54,
32'h3b1efefe,
32'h3ee789bc,
32'hbe43161b,
32'h3ddd1d9a,
32'h3ec4b17d,
32'hbedd0d73,
32'hbe7051b9,
32'h3e9e4c5f,
32'hbf5312f9,
32'h3e3823be,
32'hbf5c4b6f,
32'h3d3870a8,
32'hbc109891,
32'h3f1ac12f,
32'h3f1723e0,
32'h3f0573e6,
32'h3eadb699,
32'hbf6e1782,
32'h3e90596b,
32'hbf46d169,
32'hbe61292c,
32'h3ef73dbe,
32'h3c74b09c,
32'hbf73b01b,
32'h3ed74851,
32'h3daa3598,
32'hbf0b1c92,
32'hbf1c6554,
32'hbf5caaa7,
32'h3ecae15a,
32'h3dadd7ee,
32'h3f2beee7,
32'h3e355220,
32'h3f2eb888,
32'hbeb25d3d,
32'h3f1457d9,
32'hbed69d11,
32'h3f1642d6,
32'hbf05fc3e,
32'h3f5b6be4,
32'hbf1b744d,
32'hbd7babb8,
32'h3dec3474,
32'h3dd16193,
32'h3f963608,
32'h3f111836,
32'h3f2d7bc6,
32'hbf2916af,
32'h3ec14604,
32'hbf576028,
32'h3ee12247,
32'h3edd2c56,
32'hbed8bcef,
32'hbf852422,
32'h3ea7c356,
32'h3ecc70e5,
32'h3e6be6b2,
32'hbdb9dfcd,
32'h3c214f83,
32'h3f820997,
32'hbe0bcc3d,
32'hbf7c71d4,
32'hbe98d168,
32'h3f19aab3,
32'hbf2936a5,
32'h3f1880de,
32'hbe94f7b1,
32'h3df5fcb1,
32'h3e52094f,
32'h3f2bab49,
32'h3e364749,
32'hbc90a06f,
32'h3dc71ff3,
32'hbe6ea9e6,
32'h3f0d8a26,
32'h3dbf9bee,
32'h3eea7e99,
32'h3e8d9b7c,
32'hbae18d9a,
32'hbee390b0,
32'h3dcfdae1,
32'h3edd6c2c,
32'hbda15326,
32'hbf9136c3,
32'hbdbc1a8e,
32'h3f1a3aaa,
32'hbe0a623e,
32'h3e3d2a4d,
32'hbd3e525a,
32'h3fb1c952,
32'h3d750fe1,
32'h3d8a83b8,
32'h3d0a85b4,
32'h3ee17304,
32'h3e29a303,
32'h3d854660,
32'hbe0e2592,
32'h3d1ef216,
32'h3ea2e8dd,
32'h3ed32555,
32'h3d78b491,
32'hbca2598e,
32'hbda2bdf4,
32'h3e1b26ad,
32'h3e959e6e,
32'h3d5fed49,
32'hbe9cab7c,
32'h3e90f511,
32'hbb727337,
32'hbe3c895b,
32'hbd6ce51b,
32'hbe481d91,
32'hbd059b84,
32'hbda9f02e,
32'h3d418a1e,
32'hbde89270,
32'h3d2c3ef0,
32'h3df6cbdf,
32'h3d2e5d2d,
32'h3f2d21cc,
32'hbe0505db,
32'h3da67d28,
32'hbc506d34,
32'h3cd90f08,
32'hbd39db6f,
32'hbdca27db,
32'h3f28cfd3,
32'h3e847f8e,
32'hbcce338b,
32'h3d8f528c,
32'h3ad32534,
32'hbc236fe4,
32'h3d04af13,
32'hbd8da0ac,
32'hbd6fe039,
32'hbccdd64b,
32'hbea5c4e6,
32'h3d7123a3,
32'hbaa14094,
32'hbdb1a705,
32'hbda7ea8f,
32'h3d861720,
32'h3f059487,
32'hbd73d899,
32'h3d40f91d,
32'hbd2c8ca1,
32'hbdc9986b,
32'h3f743b68,
32'hbcbace79,
32'hbda6191e,
32'h3cbd58ec,
32'h3c9db0c4,
32'h3e139f17,
32'hbc2c276e,
32'hbd876f4b,
32'h3d60682f,
32'h3d13e01d,
32'h3f0a40ef,
32'h3e270c83,
32'hbdac523e,
32'hbbae4226,
32'h3cb744c4,
32'h3db8411f,
32'hbe1980dd,
32'hbecae663,
32'hbd49bf35,
32'hbebbfd91,
32'hbd9f3b1f,
32'hbd28b6cf,
32'h3e9634b3,
32'h3e1fc115,
32'hbd0830a6,
32'h3e0590b8,
32'hbd0313fc,
32'hbe47d3f7,
32'h3f00fa51,
32'h3e1e428e,
32'hbdec4ac3,
32'h3df7d96c,
32'hbd469ddf,
32'hbc19bf59,
32'h3ec2fca7,
32'h3f9566eb,
32'h3d97194f,
32'h3e0c872e,
32'hbd06f72f,
32'hbd74baf0,
32'hbe83e120,
32'h3f2c08ff,
32'hbe4608b5,
32'hbd2f8af3,
32'h3ca5df92,
32'hbdd3f6ff,
32'h3ec6a34a,
32'hbf59a595,
32'hbdd6ff92,
32'hbeeed04c,
32'h3f1d93f2,
32'hbed04548,
32'hbe4ef1f0,
32'hbe0e2613,
32'hbe64dd32,
32'h3f469613,
32'h3d8609ad,
32'hbeb48fe6,
32'hbf10ffdc,
32'h3f21cedf,
32'h3ef08caf,
32'h3f2e0532,
32'hbf059210,
32'hbf2fc3d2,
32'h3ea03f54,
32'h3ebc2028,
32'h3f0a4318,
32'hbf253ae9,
32'hbd9ab5eb,
32'h3d1ae89d,
32'h3e432c5c,
32'h3f43e370,
32'hbf67e2ca,
32'hbe413dda,
32'h3ccf1e9b,
32'h3d3b7ebf,
32'hbf82fe7a,
32'hbdd2ddba,
32'hbf1ffbf3,
32'h3f1e01b6,
32'h3f08f543,
32'h3e7d9166,
32'h3e1e5425,
32'hbf1c1635,
32'hbf8abd18,
32'hbf082e3a,
32'hbe922c68,
32'hbe5c6a51,
32'hbf93dac5,
32'h3f119489,
32'h3dfbf101,
32'hbcae2bf3,
32'h3f0f9465,
32'h3dc766e2,
32'hbdf0f4ed,
32'hbebd2abc,
32'hbeec9f28,
32'hbee1e727,
32'h3d26d790,
32'hbe59b166,
32'hbd2c98f0,
32'h3f2744fc,
32'hbf931cd0,
32'h3f65abe1,
32'hbd9878e9,
32'hbd48a803,
32'hbe25393f,
32'h3e74a071,
32'hbea8ad0a,
32'h3ef152d7,
32'hbe891748,
32'hbe294a72,
32'h3eef85da,
32'hbe85e6f5,
32'hbf42ef58,
32'h3ea492ae,
32'hbe61d913,
32'h3ea1ac46,
32'hbfcd77bc,
32'hbe9feb35,
32'hbe54b45a,
32'hbd463cc3,
32'hbe32cdfb,
32'h3f065a2d,
32'hbf163095,
32'hbce8201d,
32'hbf23c78e,
32'h3e4f14c4,
32'h3c36b63d,
32'hbeabff6c,
32'hbe94df77,
32'h3ee260da,
32'hbf81dcad,
32'h3dd64efa,
32'hbc8f6b45,
32'h3d2e3aca,
32'h3e6bbe7d,
32'hbf3dea12,
32'hbf7f61b4,
32'hbe86c02d,
32'hbfa13f0a,
32'h3f35a6fa,
32'h3e34f87f,
32'h3e51c792,
32'hbd22e8a2,
32'h3daa0b9b,
32'h3e835d4f,
32'h3ce80e5b,
32'hbf8014de,
32'h3ef07680,
32'hbeef6a45,
32'h3edb432d,
32'h3edffef9,
32'h3f0a464b,
32'hbec19cd9,
32'hbd26e914,
32'h3f036251,
32'h3f07d583,
32'h3df3b253,
32'hbe961bdf,
32'h3e64aff7,
32'hbebdf0ef,
32'hc001c2b5,
32'hbe8fed27,
32'hbb9607b5,
32'hbdc92a56,
32'h3e5d84aa,
32'h3e932693,
32'hbfa12b2b,
32'hbeb34238,
32'hbfcb9576,
32'h3db59c6d,
32'hbe70bdf3,
32'hbe240fa8,
32'hbbf07259,
32'h3eb788f6,
32'h3e4f331f,
32'h3e97d4cc,
32'hbfa654bf,
32'h3ccc4cb4,
32'hbe445b7b,
32'h3e0fb77c,
32'h3f501e67,
32'h3eb26a43,
32'h3eec2ac8,
32'hbe9cad6c,
32'hbdc2ecd6,
32'h3edc4f10,
32'h3e9582d8,
32'hbe3d4afc,
32'h3df0e484,
32'hbf047bff,
32'hbf993cbe,
32'hbd2861ea,
32'hbc5cf3c3,
32'hbac2b4ab,
32'h3e020396,
32'h3efca281,
32'hbf8f8f93,
32'hbe21fff8,
32'hbf6763e2,
32'h3ec0e173,
32'h3d67a415,
32'h3d979e57,
32'h3e90e9e3,
32'h3de655e4,
32'h3f014c94,
32'h3e954d27,
32'hbe3ce3f5,
32'h3e3c6330,
32'hbdf54709,
32'hbc746aaf,
32'h3f3f582f,
32'h3e5d816f,
32'h3e5e3611,
32'hbbf0c60a,
32'hbfc068fa,
32'h3ecda888,
32'hbdab5eec,
32'hbe20cffb,
32'hbc50321e,
32'hbdc8e900,
32'hbf8f1fd8,
32'h3f4a86b1,
32'hbc42acf6,
32'h3c82afca,
32'h3e9fad60,
32'h3ebc6a9c,
32'hbfd15a45,
32'hbdcb90c3,
32'hbebb01cf,
32'h3e162595,
32'hbe117198,
32'h3d2900fa,
32'h3e530200,
32'h3e5308fa,
32'h3f221c8d,
32'h3e5ce9de,
32'h3e481725,
32'h3b49165b,
32'hbd875b35,
32'h3d344903,
32'h3e838d5b,
32'h3e94c883,
32'hbed2074f,
32'h3e2282ce,
32'hc002a503,
32'h3e1b1678,
32'h3e181491,
32'hbdd72588,
32'hbe9b0599,
32'hbc18a816,
32'hbf4f6f45,
32'h3de02cdc,
32'hbcd50dea,
32'hbd5d6b93,
32'h3dda301d,
32'h3f407f77,
32'hbfb92686,
32'hbd307194,
32'hbf566f79,
32'h3ec5be18,
32'hbd7095b5,
32'h3e867b66,
32'h3e54e2b2,
32'h3e938407,
32'h3dcc74a5,
32'h3de1cde8,
32'h3e3c07e4,
32'h3d33f497,
32'hbea18018,
32'h3dec30eb,
32'h3e780b28,
32'h3ed228f1,
32'hbec29fd2,
32'h3dd5bbc1,
32'hc0068344,
32'h3e26d593,
32'hbea91eed,
32'h3e5c7109,
32'hbe84a0bf,
32'hbd88b7b0,
32'hbd38f2b6,
32'hbf6716d9,
32'hbd95d2da,
32'hbdb595b4,
32'hbd2db3e4,
32'h3dc18cd5,
32'hbfc0c46d,
32'hbae7c4a1,
32'hbe7dc786,
32'h3e9217f2,
32'h3dd3a205,
32'h3d30f1d5,
32'hbd2574de,
32'h3e136c52,
32'h3e16e055,
32'h3dd8a013,
32'h3dca8b63,
32'hbe9d0d12,
32'hbd7261fe,
32'h3e1f495e,
32'h3ec6b2cb,
32'h3ed30cb6,
32'h3ce243ec,
32'h3e9a1e3e,
32'hbefa129d,
32'h3dec2988,
32'hbe4714cf,
32'hbdebe607,
32'hbe7ad9f2,
32'hbbe439c2,
32'hbd0213f0,
32'hbeb51b8d,
32'hbca48b83,
32'h3cc2d4c2,
32'h3d465519,
32'h3e79fb16,
32'hbed4c869,
32'h3daa3201,
32'hbe0f295c,
32'h3e466d5e,
32'h3d8758ba,
32'h3db34548,
32'h3ea16e0b,
32'hbbe43850,
32'hbdc6d310,
32'h3e13d64a,
32'h3ea098a5,
32'hbf206993,
32'h3e11e45b,
32'h3e193585,
32'h3ee0d4da,
32'h3f249b64,
32'hbe3c8c3f,
32'hbe7452ab,
32'hbe1231de,
32'hbecfefc3,
32'hbea86549,
32'h3d8b3e7d,
32'hbd925e67,
32'h3db0844b,
32'hbdcea37e,
32'hbe85c312,
32'h3d9d38f4,
32'hbd8fac71,
32'h3e43e4d6,
32'h3ed51ac4,
32'hbe864bb8,
32'h3e2fb269,
32'hbe762038,
32'hbe0b4e64,
32'hbe46dd48,
32'hbd8fcca5,
32'h3e5ddf39,
32'hbcbbaa37,
32'h3ec9a09e,
32'h3e48493c,
32'h3e4f616e,
32'hbf4c3b5c,
32'h3de74fb9,
32'h3caea132,
32'h3e2d912c,
32'h3daeaf78,
32'h3e08d472,
32'hc001e786,
32'hbe1c73c1,
32'hbf481fb2,
32'hbde9ab15,
32'h3d9437da,
32'hbd93de12,
32'h3d9fa152,
32'hbd87e46b,
32'hbe9209ff,
32'hbd0b2cd0,
32'hbb974e20,
32'h3e2a28d4,
32'h3e416ac1,
32'hbf5f5fdb,
32'h3e855eff,
32'h3d154092,
32'hbe2a4870,
32'h3d9b4572,
32'hbebf0ab6,
32'h3d7381b9,
32'h3d5caf82,
32'hbdc56e0d,
32'h3d2777b8,
32'h3e3a2320,
32'hbfc53488,
32'hbd9295f3,
32'hbd2d9b2a,
32'h3de83c5f,
32'hbe9d4cf0,
32'h3e686eba,
32'hbf80ded4,
32'hbe3e2641,
32'hbf86e237,
32'h3e432f4c,
32'h3e3ba373,
32'h3eb2469d,
32'h3cab5198,
32'hbe55f90c,
32'h3ea23192,
32'hbd59eff9,
32'hbcd109fc,
32'hbd6bd420,
32'h3e3986cd,
32'hbf558469,
32'h3e871017,
32'h3dc98c0f,
32'h3dbbe1eb,
32'h3dd0762d,
32'hbf083860,
32'hbd4ce650,
32'h3cfe22a4,
32'hbea69e78,
32'hbe07b458,
32'h3eeaa802,
32'hbe75ad66,
32'hbd73fb35,
32'hbe8ce354,
32'hbd4d7a8a,
32'hbf173566,
32'hbd67aae7,
32'hbed8e64d,
32'hbe73a86c,
32'hbf810aaa,
32'h3eb33302,
32'h3d244ce9,
32'h3e8b2900,
32'hbc0578d2,
32'hbe42c5e9,
32'hbd18d881,
32'hbcb7c435,
32'hbd9e30b8,
32'hbd9103e1,
32'hbe8b1fe5,
32'hbdfe53dd,
32'h3e723608,
32'hbc551372,
32'hbd8511a7,
32'h3e05f680,
32'hbf27f175,
32'h3e6d20cf,
32'h3dfe7d28,
32'hbe926b34,
32'hbe46c115,
32'h3d5a7104,
32'h3d8c135a,
32'hbb8bc234,
32'hbd94b9df,
32'h3e2ae28f,
32'hbe94bb38,
32'h3ddce02d,
32'h3d762ece,
32'h3d18b244,
32'hbf8148da,
32'h3e6148ce,
32'h3cb11495,
32'hbe8bcb9d,
32'hbda02df1,
32'h3d7f550f,
32'h3e2d10da,
32'hbda9cbbb,
32'h3ca28b21,
32'hbea6fe3b,
32'h3ca9cc16,
32'hbed6ad42,
32'h3e419d8f,
32'h3b8847ae,
32'hbb807c8d,
32'h3e9239a9,
32'hbd919a9c,
32'h3e62db10,
32'h3e4f4dff,
32'h3da17801,
32'h3d85a69a,
32'h3e724364,
32'hbe16bb8a,
32'h3d5470ad,
32'hbe26891b,
32'h3f1a1c59,
32'h3e0870bf,
32'hbebd1829,
32'h3d22cfc1,
32'hbbedbe01,
32'hbed5819d,
32'h3d964aa2,
32'hbeabee9c,
32'hbe85e2c0,
32'h3e077a5f,
32'hbc8dd3f7,
32'hbeb14bc2,
32'hbde64600,
32'hbc5b391b,
32'hbddb7cda,
32'h3cd8cf25,
32'hbea9d215,
32'h3ebf28e1,
32'hbe69f0b0,
32'h3ec41204,
32'h3f009285,
32'h3ec6329c,
32'h3df600e3,
32'h3f02da13,
32'hbd907e9b,
32'h3d2b39d3,
32'hbd8e5508,
32'hbbd515e2,
32'h3dab59b6,
32'hbdba4726,
32'h3dd3d3a5,
32'h3e9805e8,
32'hbee9f22b,
32'hbb127c91,
32'h3e2f2e78,
32'hbe25a061,
32'h3e962614,
32'h3e050d64,
32'hbe2b0484,
32'hbe0a428b,
32'h3da94965,
32'hbf0a3a78,
32'hbd722f38,
32'h3b39f71f,
32'hbe220296,
32'hbbba648f,
32'hbdf54e5b,
32'h3e11446b,
32'h3e4e8680,
32'h3e6b59fd,
32'h3e3b4279,
32'hbdaffebe,
32'h3dacdbce,
32'h3dc83bd9,
32'hbe87df4f,
32'h3e160078,
32'h3d98e9b0,
32'hbe67d802,
32'hbe874303,
32'hbef36c3b,
32'hbe4b15fc,
32'h3d5237f1,
32'hbe8e7f67,
32'h3e859ef3,
32'h3d05b35c,
32'hbe906063,
32'h3edf6afa,
32'h3cc561d5,
32'h3c576c2a,
32'h3982b966,
32'hbc5a4145,
32'h3efa0243,
32'hbc82eccd,
32'h3da692dd,
32'h3d80d709,
32'hbe4397fa,
32'hbda5e2a7,
32'h3c988870,
32'hbf5373e2,
32'h3f0e5dca,
32'h3f01628e,
32'h3e4358cd,
32'h3ea10221,
32'hbd8b84cb,
32'h3e4fbb76,
32'hbe8c3dac,
32'hbd800c43,
32'h3e3d7bfb,
32'hbed2e933,
32'hbf70776d,
32'hbe838414,
32'h3e266159,
32'hbea61181,
32'hbe4325a5,
32'hbe1acc1c,
32'hbda66a6c,
32'h3e2c34ff,
32'hbe1a73ad,
32'hbddf16a9,
32'hbc28e44c,
32'h3d2be23f,
32'h3d9e3f61,
32'h3c41de83,
32'hba8fbaaa,
32'h3ebe161f,
32'hbe9258b6,
32'hbda8f5af,
32'h3e1c4c54,
32'hbffc4092,
32'h3e23a583,
32'h3e83c9ed,
32'hbd7cb84d,
32'h3ecc3557,
32'h3e919344,
32'h3ee398e5,
32'hbdcb519c,
32'hbd98da24,
32'hbf3c2b52,
32'h3e327fee,
32'hbfe1cc48,
32'hbdc2b0a4,
32'h3ded5cc5,
32'hbdbab5f3,
32'h3e0899ae,
32'h3e06e833,
32'h3e2151bb,
32'hbd651382,
32'hbd1bd180,
32'hbde98058,
32'hbe310fed,
32'hbe8a8887,
32'hbf0b929c,
32'h3d04e26b,
32'hbd1909a6,
32'h3e9970fe,
32'hbe9cb74e,
32'hbe8666fb,
32'hbc3e5684,
32'hbfb8487e,
32'h3e93078e,
32'h3e71aa54,
32'hbd609ae2,
32'hbc96bb0f,
32'h3e94dd38,
32'h3e9e9768,
32'hbdb0eb0c,
32'h3f142cc4,
32'hbdcb795a,
32'hbced9a5b,
32'hc01a34c4,
32'h3db879e6,
32'hbe12a5e8,
32'h3eb2c86a,
32'hbde5803c,
32'h3ddbc934,
32'h3e913930,
32'h3f0586f1,
32'h3e97640d,
32'h3d80a5c1,
32'hbbd17059,
32'hbd425f48,
32'hbef6e2c0,
32'hbd21c098,
32'h3d0c77ed,
32'h3ebda571,
32'h3de8293b,
32'hbe888b8e,
32'h3d09fc2f,
32'hbf76f138,
32'h3e6c9202,
32'h3d4e4821,
32'hbe88c699,
32'h3e6df2e2,
32'h3cf61f71,
32'h3f652767,
32'h3e89aa8b,
32'h3eb49b4b,
32'hbe1bed41,
32'hbee8ca5b,
32'hbfdb47ab,
32'hbc46387c,
32'h3ead0010,
32'hbe61821b,
32'h3f23119f,
32'hbe40a941,
32'h3e6408f6,
32'h3e1cc2aa,
32'hbecb542c,
32'h3e58ad15,
32'h3e89e505,
32'hbd48dd48,
32'hbedaedf0,
32'hbd8a3b64,
32'hbd5b839e,
32'h3ed970b1,
32'hbca3e7cd,
32'hbddf92f4,
32'hbd8bece8,
32'hbf6000a1,
32'hbe3a854c,
32'hbc6e9c07,
32'hbe3919b6,
32'h3e2407f4,
32'h3e7f9541,
32'h3d0545f7,
32'h3eb904ca,
32'h3e6d8622,
32'h3eceee09,
32'hbe7bedc9,
32'hc013c1bd,
32'h3d22dc88,
32'hbe139c3c,
32'h3f62e2d9,
32'h3f13846d,
32'hbe9afbea,
32'h3f05a06c,
32'hbee66521,
32'hbe560de0,
32'h3f4da9c1,
32'hbf0a078b,
32'h3d83e7c6,
32'hbede9fb5,
32'h3d6e6a6c,
32'h3bf034c5,
32'h3f08f4f8,
32'h3e1a645e,
32'h3e253aa5,
32'h3eb13b16,
32'hbed76a3b,
32'hbe2303fc,
32'hbf292dd6,
32'hbecef3f6,
32'hbf22f4db,
32'h3d1cb161,
32'hbf844e06,
32'h3f0ec2cb,
32'h3f45d72c,
32'hbed668ba,
32'hbee627f0,
32'hbf43edaa,
32'h3e0d42d4,
32'hbeba4796,
32'h3f6ab6fe,
32'h3f211010,
32'h3d7adb79,
32'h3ec01421,
32'h3f939005,
32'hbed59f4a,
32'h3f9c274b,
32'hbd29bc0c,
32'h3f02930e,
32'h3e33251d,
32'hbcf60bce,
32'h3c993aa5,
32'h3ea20b67,
32'hbccb3b4a,
32'hbe93f656,
32'h3ec06e3b,
32'hbe6b0556,
32'h3e2b2b07,
32'h3eb775aa,
32'h3f14efa7,
32'h3e303fe2,
32'hbefba22b,
32'hbf40720e,
32'h3e1a20d2,
32'h3edc87b1,
32'h3ee6f1f6,
32'hbf0cf382,
32'hbc95f370,
32'h3ac07713,
32'hbec46f7f,
32'hbf2e1c35,
32'h3d633be1,
32'h3f4f9598,
32'hbef0e0ed,
32'h3ef2cd85,
32'hbe9867c7,
32'h3f804612,
32'h3ef787ea,
32'h3f9013e4,
32'h3faf1852,
32'hbdade70c,
32'h3d6572d6,
32'h3e8ba786,
32'h3f2d9e3e,
32'h3e2e32b4,
32'hbd3200c5,
32'h3f6c13be,
32'h3e435d65,
32'hbf6eb2ba,
32'h3ed37ee8,
32'hbf7e1fbc,
32'hbf269035,
32'hbeea9e37,
32'hbeaf1651,
32'h3f613f3c,
32'h3d01dedb,
32'h3efe747f,
32'hbdb07a14,
32'h3f391d26,
32'hbe2124d5,
32'h3c7af6ac,
32'hbd86144c,
32'h3ef290f5,
32'hbcfbf3d1,
32'hbc836dea,
32'hbda4082a,
32'h3ed008a9,
32'h3eac1b45,
32'h3f005c7b,
32'h3e70df1e,
32'h3dc08dd6,
32'hbcf4c277,
32'h3ca961f3,
32'h3f063b3e,
32'h3de6b2c4,
32'hba406f55,
32'h3f0d8e06,
32'h3d245806,
32'h3adb05c8,
32'hbe22c76d,
32'hbe23c657,
32'hbe7234b9,
32'hbd194477,
32'hbece2150,
32'h3ee8057c,
32'h3cedf2e9,
32'h3ec33c26,
32'hbd80eca2,
32'h3f0e6189,
32'hbeb9f6c1,
32'hbc08fd84,
32'h3d0dd7c5,
32'hbd1ea2d4,
32'h3d1def82,
32'hbdc96a62,
32'h3f20e339,
32'h3e35d512,
32'h3e2dfd71,
32'h3cbd05b1,
32'h3d40b383,
32'h3d270168,
32'hbd44883e,
32'h3c9a3fef,
32'h3d786f48,
32'hbd1be212,
32'hbea8d222,
32'hbba2d708,
32'h3d8bece3,
32'hbe5c2374,
32'hbda06a57,
32'hbdbd54a8,
32'h3f1645d5,
32'h3dc0ab20,
32'h3dbb3f48,
32'hbe06f9be,
32'hbb97b6af,
32'h3f67b20d,
32'h3dc81e10,
32'h3dc336cc,
32'hbc88bbce,
32'h3d23da98,
32'hbbf6493c,
32'hbd270e65,
32'h3c8e6050,
32'h3d124866,
32'h3d3e5882,
32'hbd1ddc28,
32'hbbde97bb,
32'hbd064625,
32'hbcf34b09,
32'h3dc74847,
32'hbd9f4f77,
32'h3d082cf8,
32'hbe8c3e84,
32'hbd3a0bfb,
32'hbe7aabd2,
32'h3da539aa,
32'h3d05c231,
32'hbd49c0d1,
32'h3d473275,
32'h3c2eaf3c,
32'h3e98e5fe,
32'h3d5c1298,
32'hbcd7c9dc,
32'h3e657f3a,
32'hbd2c91d4,
32'h3dbc1788,
32'hbda26197,
32'hbca8bf6a,
32'h3d83f713,
32'h3ea4b48a,
32'h3dd8a65a,
32'h3e52649f,
32'hbdd45938,
32'hbca49f8e,
32'hbde28b26,
32'hbea3d5cd,
32'hbdb67f07,
32'h3e16d7e2,
32'hbda9d843,
32'h3b862f61,
32'h3d9c065b,
32'h3d1d573f,
32'hbe8a8629,
32'hbe732fbe,
32'hbf1595ef,
32'h3f1d854a,
32'h3ef21af4,
32'hbf73af18,
32'h3f96d376,
32'hbe217fc4,
32'hbe91a11b,
32'h3d580ade,
32'hbe34d990,
32'hbccacf7a,
32'h3f35f14f,
32'h3e201d7d,
32'h3cc9933c,
32'hbf19f7e9,
32'h3f9589cf,
32'h3e40e53c,
32'h3f166efd,
32'hbef592ba,
32'hbf6399d9,
32'h3f14e703,
32'hbdb17266,
32'h3e91f26e,
32'h3bd2d8c4,
32'hbec609d3,
32'hbe3a95ef,
32'hbd049087,
32'h3ca3222c,
32'hbee20075,
32'h3f351adc,
32'hbe106d2e,
32'h3f7d5c18,
32'h3df5f106,
32'hbe3c146e,
32'hbda421ca,
32'hbdfd655e,
32'hbe55ca12,
32'hbf6674c6,
32'hbee347d3,
32'h3dae2eea,
32'h3d2f2a44,
32'h3f8b9502,
32'h3e8cb7ca,
32'h3e7b2a8a,
32'h3da23b97,
32'h3ed73866,
32'h3ea4b24b,
32'h3e54df39,
32'h3c96270b,
32'h3c0fbdf2,
32'h3f157c0b,
32'hbf0ec192,
32'h3dd14e27,
32'h3e06f6c6,
32'hbedfec07,
32'h3f1f70ea,
32'hbcf6dd5b,
32'h3dc683a4,
32'h3df812ce,
32'h3f4eb64c,
32'hbe9d967d,
32'h3ef69096,
32'hbee4dbef,
32'h3f0e3685,
32'h3ee958fb,
32'hbd773a2c,
32'h3e7b48fc,
32'hbdb4c809,
32'hbe2d3bc5,
32'h3e3dbbfe,
32'hbf20d3e3,
32'h3ed88368,
32'hbef97eb5,
32'h3e089f06,
32'h3f4cba8e,
32'h3f0460e2,
32'hbe8b1d45,
32'hbe592ba2,
32'hbec9134a,
32'h3ed97a0f,
32'hbe02b633,
32'hbf38ef44,
32'hbee379ae,
32'h3eba16f3,
32'hbf8b4270,
32'hbeb1a42a,
32'hbcbd670b,
32'h3dbd010c,
32'h3e183773,
32'h3d35cbc2,
32'hbf6df8ae,
32'h3e136c18,
32'hbef9b418,
32'h3cea3944,
32'h3bfbacf7,
32'h3df1ac43,
32'h3def0422,
32'h3e420894,
32'hbe30e540,
32'h3e2dbccb,
32'h3d151efd,
32'h3f2f438b,
32'hbc2a66a4,
32'h3ede5106,
32'h3f5978bc,
32'h3f3b2c63,
32'hbee7d7bf,
32'h3ebd408d,
32'hbf7408ab,
32'h3ea8a6ac,
32'hbc96d453,
32'hbef52412,
32'h3d931b0c,
32'hbc14eb88,
32'hbf91925d,
32'hbf57d3ae,
32'hbd8826a7,
32'h3c81d728,
32'h3e4b5f25,
32'h3f3f845f,
32'hbe29a908,
32'hbe435668,
32'hbf6631e3,
32'h3e998c3d,
32'h3d7a6763,
32'h3e3927bf,
32'hbe3e8b52,
32'h3e6df66a,
32'h3ecf9f80,
32'h3e942fc2,
32'hbbca4d10,
32'hbdde4847,
32'h3de574e4,
32'h3ea62123,
32'h3edc8765,
32'h3e62352c,
32'hbcd84798,
32'h3e459afe,
32'hbfb0426d,
32'h3f4b9568,
32'h3e89d1b7,
32'hbf3a853b,
32'hbea84418,
32'hbe71aa04,
32'hbeff5cc7,
32'hbeb679b9,
32'hbd95fc78,
32'hbdb159d5,
32'h3eaf684c,
32'h3e0898fb,
32'hbf0f427a,
32'h3e1204f0,
32'hbe07fb81,
32'h3c648de6,
32'hbe07fcb4,
32'hbe0c00cc,
32'h3e3fdc40,
32'h3d5263a8,
32'h3eedc8cb,
32'h3e9926d9,
32'hbd841da9,
32'hbc1b1558,
32'hbd7e09ae,
32'h3ba7de89,
32'h3db7133d,
32'h3f043c29,
32'h3e985934,
32'hbcb1e592,
32'hc028560f,
32'h3e8630c8,
32'hbdb9aef2,
32'hbf133dd8,
32'hbf368b81,
32'hbf12aa75,
32'hbe9fef79,
32'h3dcb8a12,
32'hbdb039bd,
32'h3d0d684f,
32'h3ec33fa7,
32'h3ef74b6a,
32'hbe3fc134,
32'hbdc79683,
32'h3e20db3a,
32'h3dc2ab30,
32'h3e5f362f,
32'h3e65f1fe,
32'h3e6387e4,
32'h3dddd143,
32'h3ed46843,
32'h3e8a2ae5,
32'hbe1452f1,
32'hbf3204b2,
32'hbe344421,
32'h3e2452cf,
32'hbda4f332,
32'h3ef1a52b,
32'h3e74ca2b,
32'h3e894bc1,
32'hbfbbff70,
32'h3ebec8b6,
32'h3d84aad7,
32'hbe27141d,
32'hbeff263f,
32'hbe9cc292,
32'hbcdf2dcc,
32'h3f1a1c6d,
32'hbe0a0827,
32'h3da1b9fd,
32'h3e954649,
32'h3f483135,
32'h3e2320c4,
32'hbc05c73a,
32'h3f045b93,
32'h3b47f154,
32'h3ca3330e,
32'h3e06965b,
32'hbd268831,
32'hbd319a2b,
32'h3eeec4cb,
32'h3d73c2e2,
32'h3e51f71c,
32'hbf6120f9,
32'hbcdca35c,
32'h3d9cc384,
32'hbe0088e9,
32'h3edd5102,
32'hbd6779ca,
32'h3f29a23c,
32'hbee4e6bc,
32'h3e3a6532,
32'hbe509d66,
32'hbd9a1b8e,
32'hbe6cf43d,
32'hbe865167,
32'h3e0076f8,
32'hbf3c740b,
32'hbc4e4be7,
32'hbd8a2041,
32'h3dfe9ed3,
32'h3e8ca52a,
32'h3e261f8c,
32'h3d1d91cb,
32'h3ecc6af4,
32'h3e7bd7ef,
32'h3e11331b,
32'h3e81c93c,
32'hbd6ac2e5,
32'hbd8f9fc3,
32'h3ea6801d,
32'h3deec8b1,
32'h3e1fb52a,
32'hbf352fab,
32'hbe7058f5,
32'h3e6f8f6e,
32'h3d4affae,
32'h3f2b2da2,
32'h3eacc3c9,
32'h3e199746,
32'h3e1e1ed9,
32'h3e56f91d,
32'hbdf6f5df,
32'hbeb83c5e,
32'hbe14538e,
32'hbee1c08f,
32'h3e098cdc,
32'h3e704d49,
32'hbc888500,
32'h3d236e56,
32'h3eb1e8ab,
32'h3dfcc951,
32'h3f160968,
32'h3cbe012f,
32'h3dea88e5,
32'hbccd08d5,
32'h3dc4d3c5,
32'h3dda5e5c,
32'h3decf4ad,
32'hbdd06b28,
32'h3d43d674,
32'hbe03c904,
32'h3e45425b,
32'hbf2a698a,
32'h3d535d27,
32'h3bca3efd,
32'h3caf70bb,
32'h3eb9bfd4,
32'h3e4ead00,
32'hc0101d4b,
32'hbd40e736,
32'hbe051189,
32'hbdb21bae,
32'h3cbd4e62,
32'h3d3dcafc,
32'hbeb62766,
32'h3eb096ed,
32'h3e16d428,
32'hbdc273b6,
32'h3bb5eba3,
32'h3cabddfc,
32'hb9f3f454,
32'h3ed1b5ad,
32'h3a94f6cb,
32'hbdaff184,
32'hbe79992a,
32'hbea9a592,
32'h3e97ac92,
32'hbdff0216,
32'hbe87d296,
32'h3e78c5f1,
32'h3c95afac,
32'h3e94ee08,
32'hbf534e9a,
32'h3ca4577d,
32'hbe2cc80d,
32'hbe40530e,
32'h3cc44e68,
32'h3de77daa,
32'hbff4e717,
32'hbe68df31,
32'hbf03dc4e,
32'hbe215d2e,
32'h3dd7e4c4,
32'h3e757810,
32'hbeac4722,
32'h3e945892,
32'h3e32783c,
32'hbb7078bd,
32'hbcadd5ad,
32'hbec9e219,
32'h3d9602db,
32'h3e49bc82,
32'h3e61b158,
32'h3d9d22e7,
32'h3ac2b308,
32'hbe9c84dd,
32'h3c38702b,
32'h3da8b324,
32'hbd314f19,
32'hbdcd7fc8,
32'hbd9b2681,
32'h3e993ee3,
32'hbe3cd2a4,
32'h3e04e1e8,
32'hbd866cb9,
32'hbe7534f3,
32'hbe0ec51a,
32'hbe7b9acd,
32'hbf0b594d,
32'hbdb7ebe1,
32'hbf834d95,
32'h3e8b0d98,
32'hbd0cd50e,
32'h3ead7d32,
32'hbe65fe50,
32'h3cab69a1,
32'h3d884d23,
32'h3d972663,
32'hbca7c4b2,
32'hbdb9fb08,
32'h3e1bc15b,
32'h3c692b49,
32'h3eb1e3a2,
32'hbe0e3198,
32'hbd8fe3d7,
32'h3db56e9c,
32'hbeadafb9,
32'h3e26a08d,
32'h3e5fa463,
32'hbefd8b0f,
32'h3d9edce5,
32'h3ca11026,
32'h3dcd7350,
32'h3e5e601b,
32'hbdd32d53,
32'hbe80bbe9,
32'h3d3cd227,
32'hbe552338,
32'h3dc45a83,
32'hbc9023a3,
32'hbf7f6dc6,
32'h3e6f202b,
32'hbd98e162,
32'h3d5265af,
32'hbea772ba,
32'hbc9f628b,
32'hbebc9a40,
32'hbc9b031e,
32'h3d6d872a,
32'hbe031283,
32'hbe7c195d,
32'hbe34ad22,
32'h3e91e4dc,
32'hbe57cab0,
32'hbdedc4c2,
32'h3e9434b4,
32'hbee8f1f3,
32'h3f05f2ac,
32'h3ea4f1b8,
32'hbe4f4094,
32'h3bca5889,
32'h3dc83ac0,
32'hbbb63681,
32'h3e0afeac,
32'hbe183cbb,
32'h3d8d8872,
32'h3db6e305,
32'h3da94373,
32'hbe263413,
32'h3dca2b91,
32'hbebad7a5,
32'hbe79a6e5,
32'hbddae40d,
32'hbe963fb8,
32'hbe59d322,
32'h3ebce422,
32'h3eb502fd,
32'hbdbeb9f7,
32'hbd333660,
32'hbd646a07,
32'h3d4e84ac,
32'hba022346,
32'h3e051554,
32'h3eb05a7b,
32'h3ce68403,
32'h3ebb00d2,
32'h3ca020ea,
32'h3e783a7c,
32'hbd1096d2,
32'h3e44921c,
32'hbd08e42d,
32'h3c584ea6,
32'hbda8f9a6,
32'hbcbb23ad,
32'hbda8c21b,
32'h3ee1a86c,
32'h3e8256ef,
32'hbd9aa48d,
32'h3ddd6b67,
32'h3dfda0e8,
32'hbf0f1f59,
32'h3e671573,
32'hbe8c8751,
32'hbd54ac7c,
32'h3dd568c1,
32'h3e032f5b,
32'hbf1d9ed8,
32'h3d54c6c3,
32'h3d5df7d3,
32'hbe155d84,
32'h3e2dc3c7,
32'h3dd2fe5e,
32'h3db6e17b,
32'hbf0807f8,
32'h3db3de2c,
32'h3eccfe6a,
32'h3e352b69,
32'h3e5d03bc,
32'h3e0709ea,
32'h3e1cc433,
32'hbc97c0d2,
32'h3df5a12b,
32'h3ef16c65,
32'hbd7ef6e7,
32'h3d1d1f52,
32'hbc7cf8a6,
32'h3ec3ba1a,
32'hbef08a4d,
32'h3e0f956d,
32'h3dab824d,
32'hbd8c0e18,
32'h3e217291,
32'h3e7397f2,
32'hbe0bf29d,
32'h3e0f0f48,
32'hbdda1751,
32'hbf55731f,
32'hbd323e1e,
32'hbd60f372,
32'hbe75dd8a,
32'hbe80ba1e,
32'hbe1d4e23,
32'hbd058d0c,
32'hbfec0d47,
32'h3dafa7e6,
32'h3e89db22,
32'hbc92b590,
32'h3e77620b,
32'h3e225f20,
32'hbd6353d4,
32'h3dc68cb4,
32'h3e55ab89,
32'h3eadc9fc,
32'hbecf8405,
32'hbcba3b28,
32'hbe81acf1,
32'hbe674468,
32'hbf1f68e4,
32'h3e8831a5,
32'h3d83ce74,
32'hbe9d7fdf,
32'hbcbd28e9,
32'hbc6d0fa2,
32'h3d9c527d,
32'h3db6e798,
32'h3e75ac8b,
32'hbe49de6a,
32'hbd95aa6f,
32'h3ac1b131,
32'h3e9e3f63,
32'h3e47498d,
32'h3e042bda,
32'h3bfd99b0,
32'hc0199774,
32'hbca36982,
32'h3e98bc97,
32'hbb250e33,
32'h3e904f18,
32'h3d0f163b,
32'h3e8cd884,
32'h3e09f34f,
32'h3e8d500f,
32'h3f152299,
32'hbdace171,
32'hbeec5884,
32'h3c60ee06,
32'hbe1efa93,
32'hbf401f96,
32'hbd652dd2,
32'hbe8a7277,
32'hbdf0d983,
32'h3d865f47,
32'h3c017f19,
32'h3ec8c1df,
32'h3ca09679,
32'h3f173b88,
32'hbf1a7bf6,
32'h3c96507e,
32'hbc115e54,
32'h3e8a746b,
32'hbe1ebd85,
32'h3e25ff17,
32'hbbb1e166,
32'hc0121593,
32'hbe097fc2,
32'h3f1132fb,
32'h3e8b33c9,
32'h3dfe9742,
32'h3e509a9d,
32'h3ea2816f,
32'h3e4c0edf,
32'hbcb70b94,
32'h3dff3549,
32'h3e064b57,
32'hbf71447a,
32'hbd9dcb0b,
32'h3e85861a,
32'h3e88dc25,
32'h3d86b726,
32'hbc47ee8e,
32'h3e2ea0d3,
32'h3dad56e0,
32'hbe0013b5,
32'h3dc966e7,
32'hbe067df0,
32'h3e13ed4b,
32'hbe4daaa7,
32'hbd16a98a,
32'hbd7dcc50,
32'h3d56c16f,
32'h3e774f5e,
32'hbd404e8a,
32'hbea42348,
32'hbf7f3204,
32'h3cb981b6,
32'h3ef7e5b5,
32'hbd7236ac,
32'h3e9a41e2,
32'h3de99c54,
32'h3da1d400,
32'h3b39b551,
32'h3f0ec16b,
32'h3f44fde8,
32'h3c891e4a,
32'hbf8421e3,
32'hbe4db33b,
32'h3e2ee0a3,
32'h3ef5057b,
32'h3d914bb7,
32'hbe404c65,
32'h3d23ae24,
32'h3e7e6ccc,
32'h3e7c44e9,
32'h3d9f06b6,
32'h3dc66fa8,
32'h3dbbd9e8,
32'hbdefb566,
32'hbd91c81f,
32'hbd9e36bb,
32'h3e59c874,
32'hbd5d75ca,
32'hbcdbab4c,
32'hbd07d316,
32'hbf19dad7,
32'h3dd394e9,
32'h3ea2589c,
32'h3db19723,
32'h3eaf3376,
32'h3e068e3d,
32'h3f478a8e,
32'h3e8215b2,
32'h3f40d357,
32'h3ddf5e99,
32'hbeb22b79,
32'hc00729bc,
32'hbe968bf4,
32'h3ea958ce,
32'h3e56cf72,
32'hbdc9cd23,
32'hbe9cd08b,
32'h3e43a60a,
32'h3e89de28,
32'h3eee7799,
32'h3edf9a00,
32'h3e468cab,
32'h3ed98a5f,
32'hbdd548e5,
32'hbde56412,
32'h3dceaa5b,
32'h3db28f63,
32'hbea877ee,
32'hbe14cc94,
32'h3d9fcb3c,
32'hbde1a9c6,
32'hbe7e2411,
32'hbcca2394,
32'h3ce6658d,
32'h3e30bbb1,
32'hbd0dcd69,
32'hbe7d9104,
32'h3f06c5c2,
32'h3eee9d75,
32'h3ebf4582,
32'hbeafb315,
32'hbfd58b74,
32'hbe03578d,
32'h3e9d3207,
32'h3f41e99b,
32'hbf1a318f,
32'hbada4256,
32'h3f314ee8,
32'h3e41d4a7,
32'hbe285dfc,
32'h3f4791e6,
32'h3eb457e9,
32'h3ee9a24e,
32'hbc659964,
32'hbdde5d85,
32'h3c08756f,
32'h3e854fc0,
32'hbbcd3e1e,
32'h3eee07ff,
32'hbd957251,
32'h3f111469,
32'hbe593af3,
32'hbee2c129,
32'hbf07816c,
32'hbf099366,
32'h3e169151,
32'hbf645634,
32'h3f105c2b,
32'h3f625aa1,
32'hbd36bfaa,
32'h3edf25a1,
32'hbfc2b78e,
32'h3ea0bcfe,
32'hbecdf53c,
32'h3eb5052f,
32'h3ec0cfaa,
32'h3e3c1c53,
32'hbd7deb03,
32'h3e9fe737,
32'hbf298088,
32'h3fa52bc9,
32'h3e5dc396,
32'h3f210e88,
32'h3ed8e74d,
32'hbda5edb8,
32'h3dc7334b,
32'h3eef8164,
32'h3e7531b2,
32'h3e8bf5da,
32'h3e2b3119,
32'h3f075c60,
32'hbd05abc6,
32'hbf3b4aed,
32'h3e8c521d,
32'hbe90af39,
32'hbe348494,
32'hbf5ae13b,
32'h3f712e90,
32'h3e128a19,
32'h3da5f150,
32'h3e2b6574,
32'hbeba510d,
32'h3f012de5,
32'h3ddc01ff,
32'hbf484306,
32'hbd124e7c,
32'h3f3b1c78,
32'hbf8682c8,
32'h3d6f69f6,
32'hbeda90dc,
32'h3f7c690a,
32'h3efe4650,
32'h3f6d17b5,
32'h3f80d62d,
32'h3d020aeb,
32'h3d99f864,
32'h3e289b91,
32'h3f3e397e,
32'h3e5b15fd,
32'hbe8226a3,
32'h3fb4cf43,
32'hbf2190ed,
32'hbfa1ee2f,
32'h3d259f16,
32'hbeea2667,
32'hbf545009,
32'hbf7a8503,
32'h3ebf0d6d,
32'h3f37171a,
32'h3ed6554e,
32'hbe9b85dc,
32'hbdd873e2,
32'h3fa04ab3,
32'h3e767be6,
32'hbd62e09d,
32'h3c8e22a2,
32'h3f691765,
32'hbecd2646,
32'hbe0cdeb2,
32'hbdc43249,
32'h3fa21ddf,
32'h3f2e3910,
32'h3fab2cce,
32'h3de8f86d,
32'h3d368daf,
32'hbaf165ab,
32'hbea290ac,
32'h3f38105f,
32'h3da52236,
32'hbd9109ee,
32'h3f49bbca,
32'h3d11e4f6,
32'hbc75ffd8,
32'hbecc67bc,
32'hbd844cbe,
32'hbf042f93,
32'hbe594118,
32'hbfa11b7d,
32'h3ef0f57c,
32'hbafd63b0,
32'h3f98809b,
32'hbd76ee07,
32'h3f30d92a,
32'hbf4dccb1,
32'hbd130081,
32'h3d0538a2,
32'hbd98acbf,
32'h3c807816,
32'h3d0419a9,
32'hbd0492fa,
32'hbd9882ea,
32'h3da0ef2a,
32'hbd16b172,
32'h3c61e507,
32'hbba241bc,
32'hbd185bf7,
32'h3cf14a65,
32'h3c9409e1,
32'h3db2ea7e,
32'h3c9e0ac2,
32'h3cd7056d,
32'h3d53b6d9,
32'hbdb3547d,
32'hbcac49b1,
32'hbc94ab99,
32'h3e2f398e,
32'hbc356ac3,
32'h3ac301b0,
32'h3bccb6c9,
32'h3cec44ab,
32'h3db73ea3,
32'hbcce86b8,
32'h3ddcb5b6,
32'h3dd27c12,
32'h3d737605,
32'hbc2d7550,
32'hbd6ff13c,
32'hbd84dea4,
32'h3d84bcef,
32'hbca833ed,
32'h3f0544a6,
32'h3f39c3da,
32'h3dc2f174,
32'hbd8fcb01,
32'h3d69edee,
32'hbd5ac0eb,
32'hbd6fbc3d,
32'hbec26c60,
32'hbdd0459b,
32'hbe2c70b4,
32'hbd4df163,
32'hbd049ad2,
32'hbd34118d,
32'hbde4a120,
32'hbbfba02f,
32'h3e9c1d50,
32'hbcd7a11d,
32'hbf6ad66f,
32'h3f767007,
32'hbd9acaf4,
32'h3f0b7f2b,
32'hbc726c30,
32'h3e98f610,
32'h3d042115,
32'h3ec9e751,
32'h3e10cc84,
32'h3fb7f199,
32'hbeb41309,
32'hbdc6a935,
32'h3f115502,
32'h3f14b748,
32'h3eec5eea,
32'hbce8eba3,
32'hbe283504,
32'hbd4dfef0,
32'h3ca5e64c,
32'hbdea357c,
32'hbea18281,
32'h3ec65ffa,
32'hbe8dca27,
32'h3f1c7380,
32'hbdf7556a,
32'hbf8fb958,
32'h3f2fb170,
32'hbe8f2efd,
32'hbeb6f132,
32'hbd8bf8ee,
32'hbf8130f3,
32'h3f4e7efe,
32'h3efb32e6,
32'h3f554f69,
32'h3e9f8601,
32'hbef337af,
32'h3f64d509,
32'hbd82866c,
32'h3ecbee7b,
32'hbe2d305c,
32'hbfdaa800,
32'h3f0008b1,
32'h3d31cc50,
32'hbeb8bd1d,
32'hbe2f2aee,
32'h3ed5b320,
32'h3e4e8a3a,
32'hbdb425bf,
32'h3d5ae331,
32'h3ce1de68,
32'hbd91cf40,
32'hbed6072e,
32'h3f535db8,
32'hbe7499f4,
32'hbea16d4e,
32'hbf0e7da8,
32'h3da09944,
32'hbeead298,
32'h3d9b22be,
32'hbebe59fc,
32'hbe3f7459,
32'h3f5a47ba,
32'h3f1e27cd,
32'h3f342777,
32'h3e5b9f0e,
32'hbcede8cf,
32'h3e80556f,
32'hbf427342,
32'h3f6aee88,
32'hbf95b7c7,
32'h3f0459e6,
32'h3c648127,
32'hbda8a83a,
32'hbdafe9aa,
32'h3ed21b69,
32'h3e28a09b,
32'hbd8c4cd2,
32'hbdadccff,
32'h3b8a74b4,
32'h3e2d3895,
32'h3ebd9494,
32'hbf2d00b9,
32'hbd70c021,
32'h3e012a0a,
32'hbebaf387,
32'h3cade155,
32'hbea7c7fb,
32'h3e919153,
32'hbe0d66fb,
32'hbf0709b4,
32'h3d1b0f51,
32'h3f62cb03,
32'hbdf262e8,
32'hbec12f46,
32'hbcb5e68a,
32'h3f13cdda,
32'hbe9b5914,
32'hbf15669b,
32'h3cd30806,
32'hbf8d856b,
32'h3e9fb7c5,
32'h3e895b5a,
32'h3de7dd9c,
32'hbeae9c10,
32'hbd6d6a59,
32'hbe0a30de,
32'hbeb621aa,
32'hbd6fa094,
32'h3ddeb080,
32'h3dc0f4a8,
32'h3e60865f,
32'hbf26185e,
32'h3ea36415,
32'h3e7dcb7d,
32'hbe81c012,
32'hbdb7e6a0,
32'hbd90dd0d,
32'h3e266293,
32'h3daec924,
32'hbf5959e7,
32'h3e54d337,
32'h3d37f76a,
32'hbd9b68dd,
32'h3dc8bb1a,
32'h3f07fd76,
32'h3efb54b7,
32'h3e859da3,
32'hbec3052a,
32'h3ed0f64e,
32'hbfcab83d,
32'h3eef0d4c,
32'h3d57c4dc,
32'hbf07d697,
32'hbef243a2,
32'hbd161aaf,
32'h3ea9b28f,
32'h3f3deb16,
32'hbcdd461a,
32'h3d08e381,
32'h3edfae72,
32'h3f0b53a3,
32'h3e99badd,
32'h3e81c8cf,
32'h3f2b2937,
32'h3dbcbdf8,
32'h3db08294,
32'h3e4715df,
32'hbe3afcda,
32'hbdfe7cb2,
32'h3d9e0f9a,
32'h3e9120d5,
32'h3e2f35c0,
32'hbb201ad3,
32'hbd8ca8c8,
32'h3e83d293,
32'h3df7471b,
32'h3eb91956,
32'hbd2421f4,
32'h3eff9a3f,
32'hc00aca7d,
32'h3f30fe99,
32'h3e1bc527,
32'hbf54a1e4,
32'hbef2e7d1,
32'hbee93379,
32'h3e03dea8,
32'h3d903365,
32'hbd45cf72,
32'hbc4eb299,
32'h3dbfd540,
32'h3dfa0c25,
32'h3e1a1201,
32'h3e7e10d0,
32'h3f1f9468,
32'h3e600ad3,
32'h3ec5f750,
32'h3e858842,
32'hbb97fc51,
32'hbd6c06af,
32'hbb11b101,
32'h3ecb3681,
32'h3e0bd31e,
32'h3e2829b6,
32'hbe0ec0c5,
32'hbdcbcfe6,
32'hb967a450,
32'h3f1181ac,
32'h3e856e9c,
32'h3ea38f27,
32'hbfb204df,
32'h3f121100,
32'h3d9bdca9,
32'hbf9c7052,
32'hbf346334,
32'hbef3a3de,
32'hbe8bc503,
32'hbf2093ec,
32'h3cc04da1,
32'h3d25e756,
32'h3e6ecf69,
32'hbdd318b4,
32'h3eafe314,
32'h3e237971,
32'h3e4dced2,
32'hbc84a6ca,
32'h3e8672a4,
32'h3ecff562,
32'h3e48597a,
32'h3e0cf951,
32'h3e46ff00,
32'h3eb444ab,
32'h3c934cb3,
32'hbe8b8622,
32'hbde08511,
32'h3d06269a,
32'hbea9644a,
32'h3ee2f574,
32'hbda759ba,
32'h3e8aadff,
32'hbdac3834,
32'h3f0853d4,
32'hbe2595d4,
32'hbf3d4975,
32'hbed7b610,
32'hbee8569e,
32'h3d6f8f15,
32'hbd000e5f,
32'hbcf720e5,
32'h3d736f37,
32'h3e451841,
32'h3ecaf132,
32'h3ead9308,
32'h3da7000e,
32'h3e0859ad,
32'h3e66adbb,
32'hbd8d4fba,
32'h3eb0782a,
32'h3db8af89,
32'hbe390679,
32'h3e8ca6b8,
32'hbd74314a,
32'h3e656406,
32'hbf445eac,
32'h3de3af1e,
32'hbbd32858,
32'hbd7b61c1,
32'h3e955dd8,
32'hbebd0531,
32'h3f4e5930,
32'h3ebde234,
32'h3f0f86d4,
32'hbe0d5962,
32'hbee1967d,
32'hbe5552c9,
32'hbf42cd07,
32'h3cd0905c,
32'hbe0dc103,
32'hbd8294f9,
32'hbcfe014a,
32'h3eecd337,
32'h3dc3b256,
32'h3ec57383,
32'hbba0320c,
32'h3db3d2a1,
32'h3ccf4a78,
32'h3e4ba965,
32'hba840dd6,
32'h3bdab384,
32'h3d91b7fd,
32'h3e887596,
32'h3e4f29ae,
32'h3d8411cc,
32'hbf0ae5f9,
32'h3e137608,
32'h3e559ca1,
32'hbe571bac,
32'h3e845a73,
32'h3e82f8b3,
32'hbf56b79f,
32'hbbe05dec,
32'h3ede7d8f,
32'hbeb1deeb,
32'hbea56d64,
32'hbf769f61,
32'hbf8c6b4c,
32'hbd9c6a83,
32'h3daebff7,
32'hbd631c4a,
32'hbd9d2a3a,
32'h3eaa9259,
32'h3d94b51d,
32'h3eb1b3c9,
32'h3e245b2e,
32'h3e07e962,
32'hbe407bb0,
32'h3d0b78b6,
32'hbe9393ab,
32'hbde76346,
32'h3e244f37,
32'h3db7890a,
32'h3e072c33,
32'h3c529f9e,
32'hbec18cf5,
32'h3ee5119e,
32'h3e513cdd,
32'hbecfcaac,
32'h3eae41db,
32'h3d66120c,
32'hc01130d4,
32'hbc64f265,
32'hbfa24247,
32'hbdef0403,
32'hbe073ac3,
32'hbe55be21,
32'hbf8f482d,
32'hbdecae63,
32'hbe1d5028,
32'hbb171f91,
32'hbd1a8ddf,
32'hbd3edd9f,
32'hbd84f699,
32'h3dc9fd76,
32'h3e51bbdb,
32'h3e42371c,
32'h3d6f8581,
32'hbe127883,
32'hbe7f19c8,
32'hbaeaf1a2,
32'h3cf6d5d1,
32'h3e322dc5,
32'h3e21aeb8,
32'h3f0b26b6,
32'h3df8db63,
32'h3e8401a3,
32'h3cd72e7b,
32'hbec67143,
32'h3eaddbbd,
32'h3d2b5617,
32'hbf9ce3ff,
32'hbe089077,
32'hbf832c72,
32'h3e978bb2,
32'hbe12dae2,
32'h3e6b5671,
32'hbf0a599d,
32'hbb8dbf03,
32'h3dafad0b,
32'hbd43fe30,
32'h3bed9d3d,
32'hbe99d488,
32'h3d056c45,
32'h3e6ac1d9,
32'h3e649749,
32'hbdfc5d4d,
32'h3baad98c,
32'hbdf5d7e8,
32'hbd2ce6a5,
32'h3ee1ce0a,
32'h3e5b3ca5,
32'h3e6d20de,
32'hbe6a9f70,
32'h3e6be144,
32'hbe0cb663,
32'h3e83528a,
32'hbe44550c,
32'h3d87c003,
32'h3e334755,
32'hbe067737,
32'h3e20c596,
32'h3da06e20,
32'hbfc31256,
32'h3e29ff9e,
32'h3e283f17,
32'hbe7a888a,
32'hbf197fc5,
32'h3ebeded1,
32'h3da6cc15,
32'hbdb135c7,
32'hbac3bb09,
32'h3de2ccc2,
32'h3d7e9773,
32'h3e42ea44,
32'h3e5978f4,
32'hbe80c113,
32'hbd55a5e2,
32'hbd2ef026,
32'hbe97228f,
32'h3e96ba68,
32'hbd0cd7b8,
32'hbebedd57,
32'hbdc3cf78,
32'h3d85bc4b,
32'hbda2844e,
32'h3e10b10b,
32'hbe5c4d09,
32'h3e22277e,
32'h3cf9df07,
32'h3da3233b,
32'hbdb809f8,
32'hbe37a900,
32'hbef0a6d5,
32'hbe2c4468,
32'hbe77a950,
32'hbe737962,
32'hbdb6a310,
32'h3eacd9e1,
32'hbc33ddbd,
32'hbbe3ab8d,
32'hbdab9ddb,
32'hbd785356,
32'hbe407d15,
32'h3c94a954,
32'h3e6c5651,
32'hbe10f427,
32'h3e1f357d,
32'h3ebe5775,
32'hbe8968bd,
32'h3eb1d16c,
32'h3ccf03a2,
32'h3e1e705d,
32'hbdb583c7,
32'h3d7d9681,
32'hbdab34fd,
32'hbb6369c0,
32'h3deb2b3a,
32'h3ecbde48,
32'h3ead521a,
32'h3e599649,
32'hbea89cb9,
32'h3db077a5,
32'hbe513641,
32'hbdaaee7c,
32'hbe074b95,
32'hbdb71a8a,
32'hbe813785,
32'h3e93d703,
32'h3e696bd2,
32'hbd118fba,
32'hbd05b64c,
32'h3e354214,
32'h3e09b37f,
32'hbccc133d,
32'h3e43dda4,
32'h3e2c6831,
32'h3d1da5da,
32'h3e189cc2,
32'h3c328693,
32'h3ea523fd,
32'h3d84d03d,
32'h3dd295fb,
32'hbdbc3cac,
32'hbdca2eee,
32'h3e1b09b2,
32'hbe1a0e58,
32'hbd18aacc,
32'h3e109c17,
32'h3ebaf9e0,
32'hbec167a2,
32'h3e85f1e5,
32'h3e69f646,
32'hbe337732,
32'h3e1a6d61,
32'h3ca5bd09,
32'hbd43df7e,
32'h3dd4ed90,
32'h3ec37a41,
32'hbf283dcb,
32'hbbd4ea48,
32'h3c0670bc,
32'h3d78598d,
32'h3de7e19e,
32'hbb2d1228,
32'hbcb5c2d3,
32'hbfcaa42c,
32'h3d190fc6,
32'h3e8b0f0a,
32'h3d9855d4,
32'h3ed69d8e,
32'h3e721cb1,
32'h3dc35346,
32'h3d81f2ed,
32'hbc0103fa,
32'h3f02700d,
32'hbea7d8d5,
32'hbe60820f,
32'h3e8aa195,
32'h3e2c053f,
32'hbd153d42,
32'hbd73799e,
32'hbd4beffa,
32'hbd72cc76,
32'hbd437ace,
32'hbc51a9dc,
32'h3e1af8d9,
32'h3de7a234,
32'h3e6035f4,
32'hbf3da2a7,
32'h3b26c398,
32'hbdb92e5d,
32'hbbb6529a,
32'hbe8965ef,
32'h3e6e7f6e,
32'h3c81eb93,
32'hc0318ed2,
32'hbe27b2b9,
32'h3dcca5b0,
32'h3c3bc396,
32'h3f060e5d,
32'h3ec5ab32,
32'h3cfbbafb,
32'h3dc1af37,
32'hbc33fd5c,
32'h3de4595e,
32'hbe833dac,
32'hbe2b3931,
32'h3dc53a49,
32'h3c7cf17f,
32'h3e1cf889,
32'hbd9ae662,
32'h3e9801d3,
32'hbe01b063,
32'hbc9ffe31,
32'hbe75d41e,
32'h3e7a832d,
32'h3e9b65ce,
32'h3eabde42,
32'hbd4be42a,
32'hbd31efe1,
32'h3d7e59ef,
32'h3e321639,
32'h3e56ebeb,
32'hbcb9a41c,
32'hbdca5082,
32'hc0168826,
32'h3c32036e,
32'h3e2a4f4f,
32'h3d869bb2,
32'h3e2a176c,
32'h3ec60ab2,
32'hbda8aeab,
32'hbd769db9,
32'h3e892a04,
32'h3e2e17c5,
32'hbd0211c2,
32'hbb9ec20a,
32'h3eb92ad5,
32'h3e6f7c3d,
32'hbc9d59b4,
32'hbe9cacee,
32'hbe54d345,
32'h3e42ef9f,
32'h3e2ad4d9,
32'h3e77b479,
32'h3ebb87b8,
32'h3da2f5db,
32'h3e9dcd4b,
32'hbe0dd53a,
32'hbd513689,
32'hbd8bbd15,
32'h3eb80015,
32'h3ca368f8,
32'hbd87188e,
32'hbe251233,
32'hbf8eec02,
32'hbed2a872,
32'h3e5a2eaf,
32'h3e2b99df,
32'h3e65a6ec,
32'h3df2a58d,
32'h3f019999,
32'h3e9e46f5,
32'h3be73048,
32'hbe345e6c,
32'hbdd8825c,
32'hbe7d3a46,
32'h3e6d4f04,
32'h3f30b243,
32'h3edadc2a,
32'hbd0f8d3a,
32'h3e7fbf34,
32'hbd8e21c9,
32'hbcb076e3,
32'h3d9d120e,
32'h3ee9c6a2,
32'h3dfdad39,
32'h3e7e081b,
32'hbe2a224c,
32'hbcc07294,
32'hbce5c338,
32'h3df2e122,
32'h3e8e038d,
32'h3e3fd6f8,
32'hbdd39c25,
32'hbe821a49,
32'h3abb9348,
32'hbe2f7a08,
32'h3e964e23,
32'h3e9838f5,
32'h3e431de6,
32'h3e487095,
32'hbce6ee27,
32'h3e81bf57,
32'h3f302b00,
32'h3be6ee92,
32'hbf823a6f,
32'h3e5635a8,
32'h3f2b6be5,
32'h3ebc1b71,
32'hbe88e337,
32'hbd3e8a84,
32'h3bd1754d,
32'h3ebc8432,
32'h3e9e2c05,
32'h3e6dc1c0,
32'h3f429922,
32'h3e545ae9,
32'hbd4bff6f,
32'hbd5e8ce1,
32'h3cd21f8a,
32'h3e177c74,
32'h3e74ef01,
32'hbd50ad7f,
32'hbdab1034,
32'hbe715bb8,
32'hbe23f6db,
32'h3d9cb79c,
32'hbcf98c58,
32'hbe2a1419,
32'h3dea77d5,
32'h3dcfebcd,
32'hbd9d786f,
32'hbde59197,
32'h3d9a3294,
32'h3de39009,
32'hbfe4cd19,
32'h3e393976,
32'h3e6e10f0,
32'hba8498e0,
32'hbf23de2a,
32'h3ea675ec,
32'h3b029034,
32'hbec5f50c,
32'hbe9fb965,
32'h3f0fc152,
32'h3ec669dd,
32'h3ef02008,
32'h3ea10f37,
32'h3d723f22,
32'h3de567bd,
32'h3d08bba1,
32'h3e4bde5a,
32'hbe7dfc74,
32'hbdff3674,
32'h3ea49e94,
32'hbef37507,
32'h3dbca8b9,
32'hbe38a077,
32'h3ecbe439,
32'h3d1b7b07,
32'hbf0e6a57,
32'h3df2affa,
32'hbde69527,
32'hbe0a374d,
32'h3df20f75,
32'hbf7e5c9b,
32'h3dbcfc89,
32'hbdb473d7,
32'h3e5239c1,
32'hbf385ae3,
32'h3eeba156,
32'h3d311b30,
32'hbeba506c,
32'h3ea4342b,
32'h3f427444,
32'h3ad02712,
32'h3e388c22,
32'h3f8996cc,
32'h3d835f4e,
32'h3d9a1639,
32'hbdec7536,
32'hbe90c587,
32'h3e700ecb,
32'hbdb59f68,
32'hbeaf0235,
32'h3e8bd2db,
32'hbee30e5a,
32'hbde300db,
32'h3eda17b0,
32'h3e02157f,
32'h3e65d76f,
32'h3e2d0efc,
32'h3e1d7de2,
32'hbf839817,
32'h3f182817,
32'hbe9f42e8,
32'h3dae72e9,
32'h3e487a10,
32'hbe91482c,
32'hbf20085c,
32'h3fa0bcc8,
32'h3e59a8d6,
32'hbef9c524,
32'hbf97f720,
32'h3f97ca6b,
32'h3da776d0,
32'h3f81c3e1,
32'h3f8abedf,
32'hbb2c0316,
32'hbd73d2a4,
32'h3ee9bba9,
32'h3ec0f8e4,
32'h3f4054f3,
32'hbec4c7a0,
32'h3f38a598,
32'h3eb69bed,
32'hbfed9273,
32'h3e0819e8,
32'hbf17d74a,
32'hbec4b893,
32'hbf656dcf,
32'h3f4043fd,
32'h3f93ed1e,
32'hbf0bd939,
32'hbd2198d3,
32'hbeaff25c,
32'h3f1cbb0c,
32'h3e3c1b19,
32'h3ebdc7b7,
32'hbe04b08a,
32'h3f8f5b10,
32'hbfa77fb8,
32'h3f697fa3,
32'hbe758abd,
32'h3f42f42c,
32'h3e07db17,
32'h3f58bdaf,
32'h3f258511,
32'hbbcdd3b1,
32'h3df8256c,
32'hbd985666,
32'h3e8e5aa1,
32'h3e949c4e,
32'hbe07b41c,
32'h3fc9b689,
32'hbe3cff8b,
32'hbf568922,
32'h3ea5e205,
32'hbec18964,
32'hbeb3ffc3,
32'hbf6de771,
32'h3ea4836d,
32'h3e98aa18,
32'h3f339027,
32'h3d8d4d89,
32'hbe92a795,
32'h3f42fdb6,
32'hbe9d43f2,
32'hbd07e245,
32'h3dc81f27,
32'h3f592ac8,
32'hbf11277f,
32'hbe37328d,
32'hbdc9fffc,
32'h3fc4618a,
32'h3f2d9d23,
32'h3fa92442,
32'h3e19297c,
32'hbce39205,
32'hbd849af6,
32'hbe001965,
32'h3fa089cf,
32'h3d66dee6,
32'hbedf612e,
32'h3f4b292f,
32'h3d04f816,
32'hbed81220,
32'hbf082c35,
32'hbdec2736,
32'hbecfb0d8,
32'hbd74becd,
32'hbf7065c0,
32'h3f8239c0,
32'hbd2734c7,
32'h3fa1b464,
32'hbe19eadb,
32'h3f2863f8,
32'hbf94e2ea,
32'h3d64ef55,
32'hbc861a87,
32'h3d9601ee,
32'h3dac7230,
32'hbd3c51d8,
32'h3d65a2cb,
32'h3d5528f4,
32'h3dcd6d31,
32'hbbefc8fb,
32'hbde4ce74,
32'hbc3be3e9,
32'hbdc20428,
32'hbd8bbac5,
32'h3c286e5a,
32'h3ca68cb1,
32'h3c7e0157,
32'hbba2b61f,
32'h3ca5dac6,
32'hbc8fee89,
32'hbcd6f810,
32'hb9e3064b,
32'h3d87fb14,
32'hbd10aa2c,
32'hbd08e90e,
32'hbd5b213a,
32'h3db8b8ea,
32'hbdcac8b0,
32'hbd627215,
32'h3d935cdc,
32'h3d7e44a2,
32'h3e00bc4d,
32'h3b212fda,
32'hbdd16142,
32'hbd184335,
32'hbdbe8648,
32'hbd07a41a,
32'h3ee5e369,
32'h3e8c39c0,
32'h3e1c707d,
32'h3b7acd25,
32'h3d7c42ac,
32'hbd38509d,
32'hbe9d9c0d,
32'hbe64062a,
32'hbb48d17d,
32'hbf0a83c2,
32'h3d440693,
32'h3cf18367,
32'hbee9e04d,
32'h3deedf3b,
32'hbd6f4210,
32'h3e7f2da0,
32'h3c2459b6,
32'hbf5038fb,
32'h3f5fbfc4,
32'hbe1c20a8,
32'h3f22bece,
32'hbd3605bb,
32'h3eb65dde,
32'hbca87f35,
32'h3e13c0cb,
32'h3e9f51ca,
32'h3fa4735e,
32'hbee10b24,
32'hbe610a9f,
32'hbe0751ba,
32'h3ed8d2b8,
32'h3eda4773,
32'hbe3ec6e5,
32'hbc166d3f,
32'h3ca3261d,
32'h3d6242c0,
32'h3e3da581,
32'hbe0f6f1f,
32'h3ec4e47b,
32'hbda8757b,
32'hbebe4e3a,
32'hbe147842,
32'hbf888917,
32'h3f63a636,
32'h3cd4fee2,
32'hbe9063f7,
32'h3dc9385e,
32'hbf495277,
32'h3f613182,
32'h3eb87c40,
32'h3dae0f74,
32'h3eb09feb,
32'hbf002222,
32'h3f9fb94f,
32'h3f170266,
32'h3eb57cee,
32'h3ebc57af,
32'hbf896eb3,
32'h3ead5f14,
32'hbe32e4bb,
32'hbe3eeb23,
32'h3eb4ff51,
32'h3f4f0ffa,
32'h3d21dd70,
32'hbe0cc67e,
32'hbd84e90c,
32'h3d0725b3,
32'h3c02f1ed,
32'hbb90a3ea,
32'h3f003d73,
32'h3e2e87f9,
32'hbeb2e51b,
32'hbfb5192e,
32'h3e3e94ed,
32'hbebf3a40,
32'h3e784c22,
32'hbe8e7a9d,
32'hbee36dd9,
32'h3eedc88f,
32'h3e9f1431,
32'h3ef1e5be,
32'h3ed5fad2,
32'h3dd07c48,
32'hbe8cd8ae,
32'h3eb1be8b,
32'h3e917a0d,
32'hbfa5856e,
32'h3ecfde07,
32'h3eea0fb2,
32'h3dcf9ac1,
32'hbf2dd3cf,
32'h3e8fe459,
32'h3eb342d7,
32'hbc532c5a,
32'hbce36887,
32'h3cf38cb5,
32'h3cae9203,
32'h3e638781,
32'h3c8e1c01,
32'hbd092694,
32'h3dbc43ec,
32'h3e2179fe,
32'hbd0cf710,
32'h3e70e0ed,
32'h3eab3ba7,
32'hbe9373c6,
32'hbf34a784,
32'h3d213c27,
32'h3ce8102b,
32'h3e348d62,
32'hbdb8c154,
32'h3e14cab9,
32'h3da72540,
32'hbeed1be5,
32'hbeac2162,
32'hbda05e91,
32'hbf80d5f8,
32'h3d84a52f,
32'h3f17233f,
32'h3e85b927,
32'hbe975a32,
32'h3e518af8,
32'h3e740dc3,
32'h3f82198b,
32'h3c83aa65,
32'h3bfae5a1,
32'h3c9181ac,
32'h3dfebea3,
32'h3dc84349,
32'h3e97c2f2,
32'hbd44a411,
32'hbe6558ed,
32'hbd99737f,
32'hbda8989b,
32'hbebe886a,
32'h3f0194ac,
32'hbe40f85b,
32'h3f1ff3e2,
32'h3dd86d69,
32'hbe69fe96,
32'h3e260cbb,
32'h3f43b9f0,
32'h3e59f8ef,
32'hbe7ffc7b,
32'hbeac348b,
32'hbede8c54,
32'hbf8cb1b8,
32'h3e5c58c2,
32'h3e126d96,
32'h3e61fc62,
32'hbeabedc3,
32'h3e7e3433,
32'h3f549849,
32'hbe83e889,
32'hbc580a72,
32'h3c111d06,
32'h3e1bf997,
32'h3f089205,
32'h3eb819dd,
32'h3eb3fef7,
32'h3cddb983,
32'hbd857c23,
32'h3c22b876,
32'h3dd36fc7,
32'h3deb8b5a,
32'h3d6698aa,
32'hbf3665c8,
32'h3e10bd2e,
32'hbeb8840e,
32'hbf88ee0e,
32'h3db3253c,
32'h3e36e23d,
32'h3e9bc257,
32'h3e65ac3f,
32'hbe32908a,
32'h3e5f070f,
32'hbf25e472,
32'h3ec105e5,
32'hbe43f2c1,
32'hbdbe53f0,
32'hbe6ad79f,
32'h3e347d2b,
32'hbe434cc1,
32'h3d3c7119,
32'h3d323884,
32'hbdb66f5f,
32'h3db4d9ef,
32'hbe2cebd1,
32'hbd3f3973,
32'h3e62cb9d,
32'hbea22f7b,
32'h3e54bdfb,
32'h3ee1098f,
32'h3eb24664,
32'hbea407a6,
32'h3e45edbd,
32'h3d57200a,
32'h3e9679d6,
32'hbe8e00d3,
32'hbf782a63,
32'h3bd9e38c,
32'hbeade234,
32'hbd6e3ec1,
32'h3ee2994b,
32'hbecbc645,
32'hbe8ae9c6,
32'hbbc151ae,
32'h3f083c64,
32'hbe667410,
32'hbf35b966,
32'h3dd32b9a,
32'h3dc416af,
32'hbee3e284,
32'hbdb7782f,
32'hbd724139,
32'hbc8ecf30,
32'h3d03165f,
32'h3e10a3d6,
32'h3ec03b85,
32'h3ed61c57,
32'hbdb2931a,
32'hbd844653,
32'h3ed8c355,
32'h3e8a1c09,
32'h3eb5569e,
32'h3d14d29b,
32'hbc8bfd6a,
32'h3ecf3857,
32'hbed9f721,
32'hbfb1825c,
32'h3c9231ec,
32'hbf10f729,
32'h3d9212cc,
32'h3e830d77,
32'hbe1b14c3,
32'hbe9b5987,
32'h3f089547,
32'h3f1d6048,
32'hbeb3c723,
32'hbf74d9fb,
32'hbf1ebce5,
32'hbd2dcb34,
32'h3e1033ef,
32'h3e6c7652,
32'hbdc23971,
32'hbcdbf97d,
32'h3e0e102f,
32'h3e101739,
32'h3e34e5f4,
32'h3e93f482,
32'hbc35ed4c,
32'hbe444e55,
32'h3c6b207e,
32'h3e2387c3,
32'hbd8dc8ab,
32'h3ceddb81,
32'h3dbdfd10,
32'h3e9a8057,
32'hbe08e818,
32'hbf27c2c3,
32'h3d8db3f6,
32'hbe49ffef,
32'h3e523f1e,
32'h3e74592c,
32'h3d15ca99,
32'hbdf9cc14,
32'h3eb029cb,
32'h3f275ba6,
32'h3e5d7cc0,
32'hbf696ae0,
32'hbf8801cc,
32'hbd416edb,
32'h3e4ed806,
32'hbeaa12cc,
32'hbdc1cedd,
32'hbda8b56f,
32'h3e41fbf4,
32'h3e976669,
32'h3d887fb0,
32'h3eb422b5,
32'hbd6ab57f,
32'hbd93674f,
32'h3e90a411,
32'h3da3a89b,
32'h3d6a82c1,
32'h3c5ee230,
32'h3eeb0442,
32'h3e25e6d6,
32'hbe30f21d,
32'h3ef9e60c,
32'hbd5bf79a,
32'h3e1b0fae,
32'h3e249163,
32'h3f0fe52b,
32'h3e804b11,
32'hbfb068c9,
32'h3e85a80d,
32'hbe6c5f33,
32'hbda95b53,
32'hbf6eef41,
32'hbfbf2ff4,
32'hbea37243,
32'h3e094161,
32'hbe92fd2d,
32'hbd9279e7,
32'h3c49126b,
32'h3e97bb8f,
32'h3dec7abc,
32'h3e0530e8,
32'h3c4a2ed3,
32'h3d1f8a4a,
32'h3bdc5f54,
32'hbc99cf09,
32'hbe9025d3,
32'hbeb64c19,
32'h3c856784,
32'h3e16eb6c,
32'h3dfd771d,
32'hbde01ef8,
32'h3e1d3772,
32'h3e6d9b4f,
32'h3e724205,
32'h3dbb8f1a,
32'h3df851a4,
32'h3ed6fec0,
32'hbff25634,
32'h3d9dc6d6,
32'hbf8a6495,
32'h3de488a5,
32'hbece1018,
32'hbfc771eb,
32'hbef04107,
32'h3d5eee40,
32'hbda87c19,
32'hbc330712,
32'hbd0bacb0,
32'h3e1c37ba,
32'h3e511efd,
32'h3dccec4f,
32'h3e1e4c70,
32'h3df3ac71,
32'h3d077c44,
32'hbe75dbca,
32'h3d1aacd9,
32'hbe827742,
32'h3d7afcbb,
32'h3ed81c2a,
32'h3e8e1a65,
32'h3e3dc41c,
32'hbe9c0d26,
32'h3f05e969,
32'h3ddab2c8,
32'h3d2f5503,
32'hbef27c60,
32'h3e135b72,
32'hbef76d17,
32'h3e231636,
32'hbf5fbb7f,
32'h3e93286c,
32'hbebb1f71,
32'hbf6e68c1,
32'hbeefc171,
32'h3e02d47c,
32'h3eb24e41,
32'hbd9e67af,
32'h3c909c1b,
32'hbc8899f8,
32'h3ea6189f,
32'hbe23aeb1,
32'h3ee437d4,
32'hbd3da70c,
32'h3e2d57e5,
32'hbe6230ea,
32'h3e116369,
32'h3e0a001b,
32'h3e8d5b9a,
32'h3dd3a271,
32'hbe598f3b,
32'h3ea12b6f,
32'h3e045531,
32'h3e9bb9bf,
32'hbe306885,
32'h3e7d40e4,
32'h3e65d35b,
32'h3d8a4a06,
32'h3e9f7ba2,
32'h3eac606f,
32'hbf5ff3fd,
32'h3c06eaf7,
32'h3d1b74c7,
32'hbf577783,
32'hbeed3393,
32'h3d898ab9,
32'h3f01039b,
32'h3ca8e9d1,
32'hbd709d33,
32'h3e3f2cae,
32'h3ec8f064,
32'hbe80dbdc,
32'h3ed17a73,
32'hbd51ff46,
32'h3daad48e,
32'h3e037390,
32'h3e355ab7,
32'h3d030cbd,
32'h3dd2ec43,
32'hbcfe9f4b,
32'hbd835536,
32'h3e5c78ac,
32'h3d84d7e0,
32'hbe113d81,
32'hbecd4734,
32'h3e1f461c,
32'h3e893703,
32'h3d9dca76,
32'hbe71ab33,
32'h3dc01a94,
32'hbee63283,
32'h3da6aa50,
32'hbe4d3478,
32'hbeadec50,
32'hbe41d750,
32'h3da6ab94,
32'h3e277373,
32'h3d21f308,
32'h3d08660d,
32'hbd8331f8,
32'h3d6814d9,
32'hbe3dc155,
32'h3eca668d,
32'hbf25188b,
32'h3d994941,
32'h3e94fe3d,
32'h3d9fa3cf,
32'hbd368f3b,
32'h3e859f55,
32'h3e20af5b,
32'h3c0cf53f,
32'h3e7726c8,
32'hbd3da72a,
32'hbe923382,
32'h3cf04ab9,
32'h3ddac89e,
32'h3ed8a177,
32'hbf09862a,
32'hbd61617d,
32'h3bfe0aa8,
32'hbd37febf,
32'hbc7cff01,
32'hbe2342ea,
32'hbd073a80,
32'h3d382ec3,
32'hbddd73ac,
32'hbd90c6d4,
32'h3cb93540,
32'hbd2c35bb,
32'h3e0aa126,
32'h3dd64e3c,
32'h3e0c8dda,
32'h3e4ce2af,
32'hbf8690ec,
32'h3e9de4dc,
32'h3e209cbe,
32'h3e1222f0,
32'h3e86ee2c,
32'h3e2106c0,
32'h3e98c40b,
32'h3dab3dd4,
32'hbb89fda4,
32'h3e4ad3bf,
32'hbe9b74f6,
32'h3be2bd31,
32'h3da0d007,
32'h3e7be495,
32'hbed7a24e,
32'h3caf9020,
32'hbe0bdb79,
32'hbd9b8b71,
32'h3dbbee4d,
32'h3d5f1310,
32'h3da3a55e,
32'h3dad2b43,
32'hbcd637b9,
32'hbf46d6c5,
32'hbdd59e82,
32'hbd7f6e17,
32'h3ecbc436,
32'hbd4b255e,
32'h3db9bdf1,
32'hbd37a612,
32'hc0050063,
32'h3cdbf64c,
32'hbc477994,
32'h3efab88e,
32'h3e05ba57,
32'h3ed18306,
32'hbd00f31f,
32'h3d62f447,
32'hbd090557,
32'hbe1e20dd,
32'hbe7d7bbe,
32'hbe1975f3,
32'h3d9f8091,
32'h3e20b813,
32'h3eea99bf,
32'h3d3dfa90,
32'h3b16cb3d,
32'h3da2de87,
32'h3d4b57de,
32'h3e9879f9,
32'h3e59aae7,
32'hbe2e203f,
32'h3de3b6d1,
32'hbed066c9,
32'h3ca219fe,
32'hbd58e77d,
32'h3ea9d610,
32'h3d225dd6,
32'h3d31b0f7,
32'hbdabbfd6,
32'hbfb3bbd7,
32'hbd15398e,
32'h3e3fb277,
32'h3e6a425f,
32'hbdd43ff4,
32'h3e904453,
32'h3d9f6289,
32'h3bfb4498,
32'h3e01a401,
32'h3ec607fd,
32'hbe06eee3,
32'h3e39d283,
32'h3e5be662,
32'h3e12f3a7,
32'h3e62aaeb,
32'h3d961752,
32'hbdac8a70,
32'h3dbf2fe5,
32'hbe1fcff1,
32'h3df61d65,
32'h3ecc3b0c,
32'h3db39b54,
32'h3e91a213,
32'h3eb7591d,
32'h3c9b23bf,
32'hbdc0dd3f,
32'h3db1d64f,
32'hbd578ee6,
32'hbe49d6de,
32'hbd48ed01,
32'hbd274da5,
32'h3e543546,
32'hbde65d96,
32'h3ee0ac65,
32'h3d420a70,
32'h3f00b111,
32'h3ea878ab,
32'h3b4453e7,
32'hbdd8bb9d,
32'hbd047a13,
32'h3c051c60,
32'hbdb6bd11,
32'h3e72be14,
32'h3effb25c,
32'hbd95647c,
32'h3e22050f,
32'hbe6c9246,
32'h3ea17ad6,
32'h3c9ce52d,
32'h3e891810,
32'h3e2882c8,
32'hbe317299,
32'h3e9d3055,
32'h3eb19603,
32'h3cd5c6a8,
32'h3c56890e,
32'h3e8d3bed,
32'h3e0375cd,
32'hbda6bdb4,
32'hbd59103c,
32'h3f09128a,
32'hbef2d041,
32'hbcabfe79,
32'h3f02de30,
32'h3f06e56d,
32'h3f1456cf,
32'h3e270fc2,
32'h3e3c494b,
32'h3d231d28,
32'hbe8cbf2d,
32'h3d2e2ce7,
32'h3ccfe9d7,
32'hbd2d4c7a,
32'h3f066530,
32'hbdeb66b3,
32'h3eac2dc6,
32'hbe876b29,
32'hbd43f0de,
32'h3e9a9b04,
32'h3d369283,
32'h3eb3ebf4,
32'h3eeb912c,
32'hbd6f501d,
32'h3affa585,
32'h3d4311e0,
32'h3d1fed37,
32'h3e0fee00,
32'hbe9dd054,
32'h3ea38707,
32'hbe13d997,
32'h3eedad57,
32'h3e4286a1,
32'hbe5cea55,
32'h3e64d06d,
32'h3ef1143a,
32'h3ea37b67,
32'h3e47aa82,
32'h3d89c57a,
32'hbd99f5ea,
32'h3de53b57,
32'hba8e2919,
32'hbeeac3c2,
32'h3ca20067,
32'h3f128db9,
32'h3df3eb8f,
32'h3e7d9a1c,
32'hbea30889,
32'h3d704a89,
32'h3e2c4081,
32'hbbd24f2b,
32'h3e8c274e,
32'h3e0dc757,
32'hbedb88fe,
32'hbe7b9dba,
32'h3d1d8608,
32'hbc3f5a67,
32'h3eec2f1a,
32'h3b2911d8,
32'h3e157691,
32'hbd80bf3c,
32'h3e519b75,
32'hbe84670d,
32'hbe10840b,
32'hbdc44c93,
32'h3f18bc0f,
32'h3e07a788,
32'h3daf8075,
32'hbe257c54,
32'hbec31566,
32'hbe950eea,
32'h3dcb6f7d,
32'hbf90e34d,
32'h3df5e08b,
32'h3eb8b30c,
32'hbd3ecf89,
32'h3c08c6a3,
32'hbe5cdda1,
32'h3d597072,
32'h3dbdf9cb,
32'hbdd6c2bc,
32'h3ea40d08,
32'hbe4f3420,
32'h3d219b20,
32'hbe3f6904,
32'hbcfa84db,
32'hbdebca89,
32'h3e684111,
32'h3e5b9e5d,
32'h3d0733db,
32'h3d9c99d2,
32'h3eae0135,
32'hbef879ec,
32'hbe88a7a6,
32'h3edc1a05,
32'h3f14ff68,
32'h3dc7af73,
32'hbf263a93,
32'hbe59e131,
32'hbee8bece,
32'hbec5818d,
32'hbe703df5,
32'hbf8dd4d5,
32'h3edf2a95,
32'h3eca5ded,
32'h3f284fe9,
32'hbea2f89a,
32'h3ebb6d5b,
32'hbe11edc9,
32'h3e0b2aa7,
32'h3f153131,
32'h3e12efe0,
32'hbe5d1fcb,
32'h3da5230f,
32'hbf006220,
32'h3c757c79,
32'h3cd9f81c,
32'h3dc7bb78,
32'h3de321a8,
32'hbeb3de1c,
32'h3dc63533,
32'hbeec53da,
32'hbe8f50a8,
32'hbeed34d0,
32'h3e6d1aa5,
32'h3ee5475d,
32'h3e5b0899,
32'h3e4b01e0,
32'h3bb77fa5,
32'h3e401fcf,
32'h3d899695,
32'h3efe5ac2,
32'hbefa2b4b,
32'h3e76d32f,
32'h3f307875,
32'h3f31a219,
32'hbf0a9f28,
32'h3f5d6f62,
32'hbf14be88,
32'h3f5a4971,
32'hbfa7c079,
32'h3eced376,
32'h3f01ee23,
32'h3f295bfa,
32'hbc9e8cd6,
32'hbdbb9344,
32'h3c172e8f,
32'h3f3d8a0d,
32'h3f1e0f57,
32'h3fab0b58,
32'hbdd9c10e,
32'h3ec09dce,
32'h3f015a64,
32'hbf8d5395,
32'h3f423b59,
32'h3f671e1b,
32'hbed2fa61,
32'hbf18331f,
32'h3dcc666b,
32'h3f6ad1eb,
32'h3ea3a927,
32'h3d8661f5,
32'hbf28c532,
32'h3f38e226,
32'hbe43616f,
32'h3e9e739a,
32'hbe1ee9f9,
32'h3f594723,
32'hbfbd2cfd,
32'h3f0caf05,
32'hbf8f6c88,
32'h3ede3f84,
32'h3dfca5fc,
32'h3f3bbc12,
32'h3ea6d321,
32'hbda50c0a,
32'h3ccdf598,
32'hbea2b183,
32'h3f90e3a6,
32'h3f76ade7,
32'hbe92da6e,
32'h3fa5a851,
32'h3e03219d,
32'hbfaf918c,
32'h3f46c28d,
32'h3f10b903,
32'hbf03e80e,
32'hbf78aa7c,
32'h3e0e343d,
32'h3f245b0b,
32'h3e0264fe,
32'hbe395314,
32'hbef2751f,
32'h3f012b58,
32'hbf02c0ed,
32'h3ca5b6bf,
32'h3d040451,
32'h3f31aeef,
32'hbf5c4301,
32'hbdf29747,
32'hbe32885e,
32'h3fc81395,
32'h3f240426,
32'h3f82387e,
32'h3f05f224,
32'hbd8e032d,
32'h3b9fc59c,
32'hbda2859a,
32'h3f97f57c,
32'h3e1d6407,
32'hbf45102e,
32'h3fc41580,
32'h3b18659a,
32'hbeea851d,
32'hbf1bdbdb,
32'hbe490b04,
32'hbec7d875,
32'h3df1cb36,
32'hbf81630e,
32'h3f86011a,
32'hbcd411fe,
32'h3fc7a06d,
32'hbedd6c45,
32'h3f140225,
32'hbf967308,
32'hbd7d96ce,
32'h3f1f2701,
32'h3d02055e,
32'h3cfe4730,
32'h3d992868,
32'hbb89f63b,
32'h3f5636d6,
32'h3ece8251,
32'hbc8f07cd,
32'h3d22ceef,
32'hbd3be8ca,
32'hbcdd50dd,
32'hbd9c45e9,
32'hbd8f7db9,
32'hbcdfa5f2,
32'hbf0d537d,
32'h3dbb6cca,
32'hbe17fd6e,
32'h3f4da09c,
32'hbc112fe1,
32'hbf9a8749,
32'h3f187461,
32'hbbc2ee12,
32'hbf8123e2,
32'hbd93c323,
32'h3eb46f78,
32'h3f4bee2d,
32'h3eccfa27,
32'hbcf167a1,
32'hbf6a820f,
32'h3d0204d5,
32'hbc9fad84,
32'hbdb026a0,
32'h3aca7c41,
32'hbd90bf5a,
32'hbdb8162c,
32'h3f0c15ee,
32'hbe5b0942,
32'h3b8b2420,
32'h3d183c18,
32'hbc9e7671,
32'hbd89ddbe,
32'hbe6ce88d,
32'hbd986f35,
32'h3c9076b7,
32'hbea1c2e4,
32'h3e0743c8,
32'hbd86dd1c,
32'hbe732bf7,
32'h3d7c84ab,
32'h3d9f156d,
32'h3cbb8ee8,
32'h3c320e0f,
32'hbee52689,
32'h3edb4671,
32'hbd9b9095,
32'h3ddd57d5,
32'hbd9d8f23,
32'h3e28e860,
32'h3d2b0174,
32'h3d36e377,
32'h3ec591e9,
32'hbcf1cf85,
32'hbf318b1a,
32'hbea6c89f,
32'hbed57350,
32'hbd75f13a,
32'hbec49f27,
32'hbeed9f32,
32'hbdb8413b,
32'hbdce7d4d,
32'h3d801c44,
32'h3dc41bdc,
32'hbf09cc08,
32'hbb8c385b,
32'hbd8c91e7,
32'hbea32284,
32'h3d8561ab,
32'hbf580f33,
32'h3f36ba8b,
32'hbb2ce2b1,
32'hbe102d14,
32'hbd60617e,
32'hbed1c763,
32'h3e99935d,
32'h3ed8260d,
32'hbe797680,
32'h3e0cd048,
32'hbf3dcd23,
32'h3fbfac0d,
32'h3f1cf34e,
32'hbea0f00c,
32'hbf1e75d3,
32'hbf9441af,
32'h3eab3b7c,
32'hbf0c3577,
32'h3efd7278,
32'h3ef88efb,
32'h3e263626,
32'hbe9f6f07,
32'h3d16edc4,
32'h3d708bb7,
32'hbf13e4be,
32'hbe43cb7a,
32'h3e8df4d3,
32'h3e1557fd,
32'hbda4bdcc,
32'h3f1e79c5,
32'hc011fc51,
32'h3e905d53,
32'h3f6b7cc1,
32'h3de89302,
32'hbf04364f,
32'hbf1c5902,
32'h3f57766b,
32'hbf83c09c,
32'h3ed69fe6,
32'h3ea454d8,
32'h3e4d97f8,
32'h3f049d57,
32'hbeaec996,
32'h3eff89b0,
32'hbf023621,
32'h3c9444c3,
32'h3e954296,
32'h3f057619,
32'hbf455e3f,
32'hbdf7e5c3,
32'h3e8a0efd,
32'hbdebba75,
32'hbd0d158e,
32'h3d46f9ec,
32'h3ecd231c,
32'hbe06a15c,
32'hbcfefe55,
32'hbc9d3b21,
32'h3eeb896c,
32'h3e54f2fe,
32'hbf21672e,
32'hbd504ea1,
32'h3f0c9397,
32'h3d9f40b7,
32'hbf245c7a,
32'h3ebb9e60,
32'h3eab95df,
32'hbe431616,
32'h3edca900,
32'h3e526f5b,
32'h3ec836d2,
32'h3e82b3ea,
32'hbf93a2d4,
32'h3ea30733,
32'hbed93c1d,
32'h3e293439,
32'hbceaea21,
32'h3e9af3ee,
32'h3e780b93,
32'h3f079c13,
32'h3e8182d1,
32'h3d983b1a,
32'hbc854086,
32'h3daa5a9f,
32'hbe209b0e,
32'hbd809648,
32'hbc8cb9cc,
32'h3dbfa617,
32'hbf4322e6,
32'h3d0c62e3,
32'h3dcffd02,
32'h3dc0dc46,
32'hbe47dc8f,
32'h3e84082c,
32'hbefa52ce,
32'h3e9ea257,
32'h3c778477,
32'hbe0f07ab,
32'h3e80c356,
32'h3e5d0ed6,
32'h3ed5286b,
32'hbe9f0a9e,
32'hbf4b3bb0,
32'h3e4fb38f,
32'hbe25c9ff,
32'h3e355414,
32'hbdfe230c,
32'h3e3eca76,
32'h3f0f97fd,
32'h3e9b57b9,
32'h3e96feb7,
32'hbfacaa69,
32'hbca4293a,
32'h3c9351c3,
32'hbd1a4675,
32'h3f05ea5e,
32'h3e232518,
32'h3e0bd7e0,
32'hbebd746f,
32'h3e561419,
32'h3e30bfc5,
32'h3e91ee32,
32'hbccb105e,
32'h3e9ad3ee,
32'hbfa175ac,
32'h3e476ab5,
32'hbea48ec2,
32'hbed81cd1,
32'h3c62f73e,
32'hbdab0b1e,
32'h3db9a13b,
32'h3d9c7b80,
32'hbeefee3f,
32'h3e9a1e79,
32'h3f043780,
32'h3e9448f0,
32'h3dc96e1c,
32'h3eeddd9d,
32'h3e83bc16,
32'h3e9078fe,
32'h3d740d34,
32'hbea59fd0,
32'h3cc10c39,
32'h3d1186a4,
32'h3eac726f,
32'h3ecf1b07,
32'h3e3f700b,
32'h3e326564,
32'hbe953204,
32'h3e51ef2a,
32'h3f0c95e2,
32'h3ed00713,
32'hbeae8467,
32'hbe14fc70,
32'hbe715199,
32'h3ee6581a,
32'hbef81065,
32'h3d69a80a,
32'hbeb1c863,
32'hbee08866,
32'h3e1da564,
32'h3f062c7b,
32'hbdfadfe7,
32'h3ec59bd7,
32'hbe5f22fb,
32'h3f0e1893,
32'hbe866468,
32'h3ee3bb12,
32'h3e445d38,
32'h3f025b5d,
32'h3d664fc9,
32'h3dde410c,
32'hbd4e5507,
32'h3c518a21,
32'h3e0b782e,
32'h3ec60841,
32'h3ebfacd2,
32'h3e82c295,
32'h3e29910e,
32'hbd601c9e,
32'h3e40ca69,
32'h3e9c1588,
32'hbf104970,
32'hbc8c1d32,
32'hbd8a3f32,
32'h3f09812b,
32'hbf075a62,
32'hbe4bd9cb,
32'hbe27c90c,
32'hbf1b21e9,
32'h3e8e805b,
32'h3d823eb2,
32'h3d0de832,
32'hbe4c1338,
32'h3d4c1d76,
32'h3f2a7eb1,
32'hbf1a8b7a,
32'hbe7f1465,
32'h3d092a61,
32'h3f128bd4,
32'hbcc64052,
32'h3da6e9a2,
32'h3c4df9f8,
32'h3d1c0668,
32'h3def3b24,
32'h3e513882,
32'h3e972c92,
32'h3f330b3c,
32'h3ea9d822,
32'h3e45961a,
32'h3ea6cad6,
32'h3e9fb154,
32'hbf08250a,
32'h3e316e8a,
32'hbb1ca2c9,
32'h3ef32917,
32'hbce8831c,
32'h3e4b83ac,
32'hbe240ba4,
32'hbf14151c,
32'h3d8351cd,
32'h3e96cb3c,
32'h3e21df82,
32'hbf6c8a7e,
32'h3e38ed47,
32'h3f137379,
32'hbe26c0e2,
32'hbf1c3549,
32'hbe1b09ac,
32'h3ef67e64,
32'hbe1fe697,
32'hbdae3ec0,
32'hbc63866a,
32'h3cd2132c,
32'h3ed0304e,
32'h3d05b4bd,
32'h3e0ff965,
32'h3f5a0e8a,
32'h3eb02556,
32'hbd6bb8f3,
32'h3ec1d735,
32'hbe3bdf3e,
32'hbe541e96,
32'h3e9be71a,
32'h3e55a3c1,
32'h3f019a2f,
32'hbef6cb45,
32'h3ed94739,
32'hbddb8756,
32'hbec85ad6,
32'hbe20c4f0,
32'h3efdfee6,
32'h3ec5b1ee,
32'hbfa7a046,
32'h3ed35511,
32'hbd34e22e,
32'hbe898798,
32'hbf059363,
32'h3c26b75d,
32'h3eff20f3,
32'hbd7c51d7,
32'hbe4c4acc,
32'hbd7ab29e,
32'hbdb1165d,
32'h3eaf5e4d,
32'h3e826e26,
32'h3e58f205,
32'h3f57a35e,
32'h3f137af9,
32'hbe1cc4cc,
32'h3dd8d20a,
32'hbe8c6eed,
32'hbc2fa5c5,
32'h3e6849e0,
32'h3ed2fea9,
32'h3f2b25bd,
32'hbed078c9,
32'hbe0235f4,
32'h3dc191e5,
32'hbe6f36cb,
32'hbe4f8e18,
32'h3e08dbbb,
32'h3ec7f044,
32'hbf03ec54,
32'h3ea6c184,
32'hbf4f5c3f,
32'h3e8cbd6e,
32'hbf345e61,
32'hbe706091,
32'h3f34140a,
32'hbc82b9cc,
32'hbe843bfd,
32'hbc3fa13d,
32'hbbe14b36,
32'hbd7fc645,
32'h3e8b990b,
32'h3e854174,
32'h3f494fec,
32'h3e5d5a88,
32'hbd8afd22,
32'hbe2d91c9,
32'hbe096205,
32'h3db701f6,
32'h3ebb8adb,
32'h3f10f07e,
32'h3f2984fd,
32'hbdc272ba,
32'hbe894105,
32'h3e3f2f50,
32'h3e6d9867,
32'hbe0b456a,
32'h3eee3dac,
32'h3e6e9856,
32'h3edb0175,
32'h3ec6a551,
32'hbf1219e0,
32'h3eb20f92,
32'hbe253dfd,
32'hbf197158,
32'h3ed91913,
32'hbe9925f0,
32'h3e92f0a1,
32'hbd720053,
32'hbd9565eb,
32'h3e7fc8b5,
32'h3e9e50d9,
32'hbc3a3c5f,
32'h3f28a5ca,
32'hbe577843,
32'h3e82d12a,
32'h3e84a709,
32'h3e02e28b,
32'h3d691538,
32'h3e90d0a6,
32'hbe9bf6a1,
32'h3e860fbc,
32'hbe164d7a,
32'h3eaf6ef3,
32'h3d027f5b,
32'h3d63a710,
32'hbda666b3,
32'h3f225597,
32'h3c008658,
32'h3ef06e97,
32'h3e9db76c,
32'hbec7d2d0,
32'hbe16b144,
32'hbce04858,
32'hbf1d298e,
32'h3e2da3bb,
32'hbd96d005,
32'h3ee06b17,
32'hbe37b7d1,
32'h3ce5b5f1,
32'h3efad60c,
32'h3e78cc8d,
32'h3d5f0c3a,
32'h3e9d465f,
32'h3d154b1c,
32'h3e17343c,
32'h3eaf9105,
32'h3d83cdb8,
32'hbe489cb8,
32'h3db2e7da,
32'h3e9cd24a,
32'h3ee8fa64,
32'hbdb07292,
32'h3eda1b14,
32'hbeb41aaa,
32'hbdd7b8b1,
32'hbd8413c4,
32'h3e2137ee,
32'hbee6376b,
32'hbe12fd75,
32'h3e1eb43b,
32'h3bbbfc17,
32'hbdd046af,
32'h3d66ef24,
32'hbe3af730,
32'h3d3578c6,
32'h3c798ea9,
32'h3d62d2ee,
32'hbdf8a6c0,
32'hbd850547,
32'h3e59fe76,
32'h3dc339ee,
32'hbc0cab61,
32'h3eb66b80,
32'hbf80943f,
32'h3c98767f,
32'h3e1fe8b7,
32'hbcfef9c5,
32'hbd01215f,
32'h3e6bd224,
32'h3ea81a02,
32'h3ea9a939,
32'h3e0d3798,
32'hbe671d08,
32'hbe72cd38,
32'hbba71b32,
32'hbd90224c,
32'h3dfad619,
32'hbf3060ab,
32'h3bf2f14b,
32'h3e0488b0,
32'hbcfbd331,
32'h3e7378c1,
32'h3dc080ca,
32'h3e280a01,
32'h3cc5433c,
32'hbe62269e,
32'hbebb61b4,
32'hbd9f9406,
32'hbd871d70,
32'h3e1de0b9,
32'h3e4bdb18,
32'hbd5ad649,
32'h3d1ca9ce,
32'hbf8f7823,
32'hbe23750a,
32'h3d7dfe34,
32'h3e14512d,
32'hbe4c5a02,
32'h3e918248,
32'h3ec3cb4b,
32'hbc358171,
32'h3e66fdfe,
32'h39d13743,
32'hbdfdc8ef,
32'h3e013719,
32'hbd41fbda,
32'hbcb01573,
32'hbf0236f5,
32'h3d2f7ee4,
32'h3d819644,
32'h3e39629c,
32'hbe73be52,
32'h3dde3958,
32'h3e577127,
32'hbe03ad20,
32'hbd16b823,
32'hbe235637,
32'hbc27dca6,
32'hbd5dddcf,
32'h3edf6729,
32'hbb6f9e7c,
32'hbde83920,
32'hbc70b75f,
32'hbf5731c0,
32'hbddc64a5,
32'h3e03c853,
32'h3e0e5ffb,
32'hbf0c27a2,
32'h3de9c780,
32'hbe7df3d3,
32'h3e2cbe84,
32'h3e8d5158,
32'hbd99c32f,
32'hbe30756e,
32'h3ee356ba,
32'hbda8add2,
32'h3dbc300d,
32'h3eab75cc,
32'h3e5a9cd0,
32'h3e0732ee,
32'h3e42447a,
32'hbe46c9b5,
32'hbdfb6f53,
32'h3e359471,
32'hbe8ee803,
32'hbd88d2c3,
32'h3e8a02ea,
32'hbbb36309,
32'hbcf68a83,
32'h3e7f8051,
32'h3df6e866,
32'h3e3ddfd7,
32'hbc7cb6d2,
32'h3da9d212,
32'h3e01e84e,
32'h3d083002,
32'h3e8c132b,
32'hbe4aec38,
32'h3de2e31b,
32'h3cb8aeff,
32'h3ea16b43,
32'h3e2a1edf,
32'hbd89a2b1,
32'h3d742323,
32'h3ea04b83,
32'h3d794041,
32'h3e43d24b,
32'hbc38db86,
32'hbc6902e9,
32'h3e45ede7,
32'h3e080502,
32'hbebed063,
32'hbdf23850,
32'h3ebd917b,
32'hbe319f38,
32'h3db4cb99,
32'hbd8d7879,
32'h3d227b1f,
32'hbd3ea9f2,
32'hbde71d6e,
32'h3df1ff0b,
32'hbe2152f6,
32'hbd8d777a,
32'h3f17e9a0,
32'h3d12eb73,
32'hbde4169b,
32'h3dfebef1,
32'hbf0882e0,
32'h3eb7081c,
32'h3ee86aca,
32'h3e9f167d,
32'h3e7df159,
32'hbeca076e,
32'h3e1d7d2e,
32'hbe5eb4d2,
32'h3e334ab9,
32'h3e89d70b,
32'hbfca2188,
32'h3ecee770,
32'h3cb09ad5,
32'h3dbac39c,
32'hbeb8ed13,
32'h3d89ec52,
32'h3e9d7fda,
32'hbe1cd4fa,
32'hbe28f657,
32'h3ebc2ccb,
32'hbd0d04f2,
32'h3c3f6997,
32'hbdb143ea,
32'hbe250bb0,
32'hbe85033a,
32'hbd7606a8,
32'h3ee74e71,
32'hbd3deb60,
32'h3925b7b9,
32'h3d5b79c3,
32'hbef27a9f,
32'h3ec89425,
32'h3e491ce3,
32'h3d8f1b19,
32'hbd92e263,
32'h3e7aa63d,
32'h3e9b32ef,
32'hbcae2553,
32'hbe39df42,
32'h3dae324c,
32'hbe586810,
32'h3f294852,
32'h3e540a7c,
32'h3e37f6ea,
32'h3e54751e,
32'h3e051da6,
32'h3f7180f1,
32'hbe9a7949,
32'h3db1666a,
32'h3e824814,
32'h3c4d42dc,
32'h3c0ff2b2,
32'hbd2d3a08,
32'hbd8e7480,
32'h3e4c165c,
32'hbdd6a8d7,
32'h3f1fc633,
32'hbd1f574d,
32'h3dea89b2,
32'h3e9c7141,
32'hbeb4e72c,
32'h3e2eb38f,
32'h3e3e338e,
32'hbdb24ed3,
32'h3d9c08e2,
32'hbea74919,
32'h3dc1b36d,
32'hbe868675,
32'hb987c7f3,
32'h3e868796,
32'hbf56f0aa,
32'h3f0f72e6,
32'h3d762443,
32'h3e4265b7,
32'h3dc4d30c,
32'h3d944054,
32'h3efd2f7e,
32'hbe97611e,
32'h3e228370,
32'h3eab1ed3,
32'hbd36a9a3,
32'h3ca8170b,
32'hbe301c6a,
32'hbd341202,
32'h3d9daf74,
32'h3dcdd783,
32'h3f35becb,
32'hbf09692b,
32'hbefce3ba,
32'hbe5eea1d,
32'hbe406bb7,
32'h3e738bc2,
32'hbf500703,
32'h3d462abb,
32'h3b1e4dec,
32'hbf800f04,
32'h3e5e02cc,
32'hbe6e5dc4,
32'h3e1512f0,
32'h3e8d715d,
32'hbd9dcd62,
32'hbf2b09a8,
32'h3da3d8f0,
32'h3dee7b11,
32'hbe7f0798,
32'h3f11b50b,
32'h3d3b7065,
32'hbf3751ee,
32'h3e04a8da,
32'h3eb690d1,
32'h3dddedae,
32'h3dbbc383,
32'h3f16c497,
32'hbd732085,
32'h3d5d3da4,
32'hbe1633b1,
32'h3f03ad02,
32'h3e5cdd96,
32'hbf760952,
32'h3e084d87,
32'h3e9425f4,
32'h3e9118ea,
32'hbf67f321,
32'h3e8bffcf,
32'hbf0c0b3c,
32'hbf188d45,
32'h3ddd05d3,
32'hbf3595fb,
32'h3e54ff6f,
32'h3ec2d191,
32'h3e645fc1,
32'hbef50dc1,
32'h3ee33fb6,
32'hbdc336cf,
32'hbedae829,
32'hbdcf3200,
32'h3c879c0f,
32'h3f1e9988,
32'h3edec85a,
32'hbe272c68,
32'hbd450a46,
32'h3d98d3bd,
32'h3e6e67ed,
32'hbc99ba9c,
32'h3e2feb76,
32'hbe784eaa,
32'h3e3c14b2,
32'h3dee5aa6,
32'hbfa4a8c2,
32'hbde4cde5,
32'h3e934f1f,
32'h3ee72954,
32'hbfb503ff,
32'h3e6d7763,
32'h3e237315,
32'hbf16686f,
32'h3e8f5cae,
32'hbead321c,
32'h3f00abdd,
32'h3f23f582,
32'h3f2c8e05,
32'h3c248b53,
32'h3fa1ae53,
32'hbf3a4913,
32'h3eb6390d,
32'h3f223319,
32'h3efa72e6,
32'h3f397752,
32'h3f857789,
32'h3f334428,
32'hbd101409,
32'h3cd595ee,
32'h3ee820b8,
32'h3f6f215f,
32'h3fa21d16,
32'hbdeb53bc,
32'h3f55358a,
32'h3e59c8d3,
32'h3dbdd988,
32'h3e4cd18c,
32'h3f03d075,
32'hbfa573d3,
32'hbfbf92c0,
32'hbf564d6b,
32'h3f93f981,
32'h3e90e01b,
32'hbf029d3b,
32'hbf03e7de,
32'h3f2f46a7,
32'h3df63cca,
32'h3f124be5,
32'hb9f8db96,
32'h3f7560b3,
32'hbf7bdb03,
32'h3f68f935,
32'hbd895346,
32'h3e8a842c,
32'h3e134c34,
32'h3f3eebf2,
32'hbda997e8,
32'hbdb2adcc,
32'h3e24a816,
32'hbf9e7517,
32'h3f82850f,
32'h3ebcfd7e,
32'h3e95cbdd,
32'h3fa8eabc,
32'hbcc29409,
32'h3df0776c,
32'h3f1c3d12,
32'h3f97e114,
32'hbe2a2596,
32'hbea14494,
32'hbf1ad72c,
32'h3f7c1a81,
32'h3e61bf93,
32'hbd7ef2a0,
32'hbe011a29,
32'h3f0a5b33,
32'hbed7aeab,
32'h3f5ebce6,
32'h3dd55319,
32'h3e1cbcf6,
32'hbf197c3b,
32'hbd60430a,
32'h3edcebd5,
32'h3f7c454b,
32'hbe332274,
32'h3f0a37c1,
32'h3fa90c03,
32'hbd3fd567,
32'hbd6a6f01,
32'hbecf2573,
32'h3f8210da,
32'h3e161a50,
32'hbf4eea06,
32'h3f6801c3,
32'h3d7ab3f6,
32'hbe97a7ce,
32'hbe6e750e,
32'hbee90816,
32'hbf05eccc,
32'hbef3dd99,
32'hbfa24f77,
32'h3e925f56,
32'hbdfbbdc0,
32'h3f201ffd,
32'hbe3ebca5,
32'h3eaa7107,
32'hbf17296a,
32'h3cf1f272,
32'h3b6ae232,
32'hbd3dcc01,
32'h3d6b0373,
32'hbda03c4a,
32'hbcb7e69c,
32'h3cd3f582,
32'hbd656783,
32'h3c7814bc,
32'h3d88b661,
32'hbb8213f2,
32'hbddd0631,
32'h3d5a02f2,
32'hbc3496e7,
32'h3d0501a4,
32'h3c94fec3,
32'h3e24b22b,
32'hbd2e1250,
32'hbd19b5e9,
32'hbca16700,
32'hbdafbe4d,
32'hbe15cccc,
32'h3d1b36d8,
32'hbdfb1c35,
32'hbc7290db,
32'hbd80f656,
32'hbd807b92,
32'hbde3d454,
32'hbdb06303,
32'hbca207dc,
32'hbd4cb53b,
32'h3f57699a,
32'h3e2c1ee3,
32'h3d9fc5c7,
32'hbd108d5a,
32'hbdc29d7a,
32'hbc1049ea,
32'hbcbad0e4,
32'hbc782cf8,
32'h3e1ed28d,
32'hbdbca7fb,
32'hbd479cbd,
32'hbd72ec95,
32'hbe3f3cf8,
32'h3de8d62d,
32'hbf43bdb4,
32'hbd228984,
32'hbc428a49,
32'hbd696f55,
32'h3d4c0f25,
32'hbf546fdc,
32'h3f930298,
32'h3c082777,
32'hbe238a83,
32'hbefffd41,
32'h3e8f5be5,
32'h3eabda29,
32'h3da8eee7,
32'hbd6b18e6,
32'hbf717e72,
32'h3f0010b9,
32'h3f4ce409,
32'hbdd09819,
32'h3fc6bf02,
32'hbece99ac,
32'h3f915d33,
32'hbfaf7cc0,
32'hbeeac757,
32'hbf1c6713,
32'hbdd134f3,
32'hbcecc051,
32'hbc8c31a5,
32'hbdf9b50c,
32'hbef45176,
32'hbf137edc,
32'h3e9574a1,
32'hbf178f18,
32'hbe8bad3c,
32'h3efd7200,
32'h3f1a291f,
32'hbf236a0d,
32'h3f1c3395,
32'hbe0485c8,
32'hbebd596f,
32'hbeec3dfe,
32'h3f7691a8,
32'h3fac5dca,
32'h3ee0e1b7,
32'h3e8a1c1e,
32'h3e81c9d5,
32'h3ecc1afb,
32'hbf34b2cc,
32'hbf4efb01,
32'hbeb41771,
32'h3eec3aaa,
32'hbf33ad5f,
32'h3eb34c54,
32'h3f520135,
32'hbe3cb16a,
32'hbeb894c6,
32'hbb7c21ce,
32'hbbbb038a,
32'hbf1b07f3,
32'hbf517114,
32'hbdac5810,
32'h3e2ae4f8,
32'h3f276b9b,
32'h3f5e22be,
32'hbfd275d1,
32'h3ec134ab,
32'h3f5fc458,
32'h3ebbbf87,
32'hbed481ea,
32'hbd906746,
32'h3f057d52,
32'hbedc59f6,
32'h3e3ef144,
32'h3e16d10f,
32'h3d7104bd,
32'h3f4e8c99,
32'h3d25997f,
32'hbd8a716c,
32'hbdc13c0e,
32'hbd298712,
32'h3da6aada,
32'hbe7414b2,
32'hbe8486e1,
32'h3c8c7778,
32'h3ec826db,
32'hbdacc70a,
32'h3d3e654e,
32'h3da152cf,
32'h3e7e5745,
32'hbe413c63,
32'hbe0801c1,
32'hbd8ce848,
32'h3f3a7aed,
32'h3d77f679,
32'hbffc2f18,
32'hbdac77f2,
32'h3f5ebf1b,
32'hbd425b9c,
32'hbf58e3c2,
32'h3e439553,
32'h3e75b376,
32'hbe8b5b0e,
32'h3e0bc8a2,
32'h3f083196,
32'hbd88bc57,
32'h3e0d7c23,
32'hbf81b3e8,
32'hbe52ec26,
32'hbeb859c1,
32'h3ebcfdb2,
32'h3db23309,
32'h3e2225c0,
32'h3ead712b,
32'hbdb303a1,
32'h3eb785b6,
32'hbe4defcf,
32'hbd8a4401,
32'hbdb30ae2,
32'hbccbab5a,
32'h3d2ae244,
32'hbdcd63b7,
32'hbe9dd400,
32'h3df44387,
32'hbcd5792e,
32'hbf382efc,
32'h3e186de0,
32'hbe4e5c10,
32'hbdc9c5b5,
32'hbfa668d6,
32'h3c8d7eeb,
32'h3e95e900,
32'hbcabfc01,
32'h3ca6d192,
32'h3eda56e0,
32'h3e68c5d2,
32'hbed6a3ab,
32'hbf05f1b7,
32'hbe67cec5,
32'hbdb88e80,
32'h3e1510a1,
32'hbeff10cf,
32'h3e37d096,
32'hbb2490a0,
32'hbe0860a8,
32'hbd3f8ce7,
32'hbfa4a71e,
32'h3c43610c,
32'h3d1c0b5a,
32'hbcbad8d7,
32'h3d6ce298,
32'h3ec61418,
32'h3d20b22a,
32'hbee4fe4b,
32'h3e28f787,
32'hbe2d07ce,
32'h3ecdeb96,
32'hbedf4ed1,
32'h3e9fa9d8,
32'h3dccec01,
32'h3e157482,
32'hbde57b7a,
32'hbf2f8a2b,
32'h3e3256e2,
32'h3ed558cc,
32'hbdf6eb08,
32'hbea6f8fb,
32'h3e4a3348,
32'hbd3b40df,
32'h3e6e1921,
32'h3e85edcc,
32'hbe964753,
32'h3daa248f,
32'h3e84c535,
32'hbd06d766,
32'h3d923cc9,
32'hbea21ffc,
32'hbc9a2544,
32'hbd5f45fb,
32'h3e068058,
32'h3e73a877,
32'h3f1cc024,
32'h3e646fb5,
32'hbdcddbc5,
32'hbea048e2,
32'h3eb498fe,
32'h3e502074,
32'hbfbf1927,
32'h3dcd33b4,
32'h3e175f91,
32'h3e45b53d,
32'hbebe4d58,
32'h3e0b07da,
32'hbcecd74f,
32'h3e5f352d,
32'hbd73930c,
32'h3c8059e2,
32'h3da71c97,
32'hbf07bf47,
32'h3c7a8f21,
32'h3e8bdd57,
32'hbec0d51a,
32'h3e7b5593,
32'h3e5d669d,
32'h3dd985d3,
32'hbd8b9cca,
32'hbf069402,
32'h3c654332,
32'hbcae36e2,
32'h3e887d68,
32'h3e1be743,
32'h3e71f997,
32'h3e7c7cd6,
32'hbd498566,
32'hbdc78b32,
32'hbd67fab4,
32'h3ed536e5,
32'hbfcc0a36,
32'h3ea06d48,
32'h3da0caae,
32'h3f0e3128,
32'hbedaf7ab,
32'hbdc5b9f1,
32'hbd3c99c5,
32'h3d20b138,
32'hbe07bd76,
32'h3e3047da,
32'h3e110398,
32'hbf989d92,
32'hbc8f2dd5,
32'h3f535a19,
32'hbe08241a,
32'h3eb483bc,
32'h3e162700,
32'h3e997e13,
32'h3ca64d6a,
32'h3e922a66,
32'hbc7c5d15,
32'hbd4db46f,
32'h3e9ae6de,
32'h3e264b0f,
32'h3e62080d,
32'h3ec8dd17,
32'h3e7ee9e3,
32'hbe6df652,
32'hbd3e59b1,
32'h3e8e05b5,
32'hbf931a02,
32'hbc66c72f,
32'h3ec09130,
32'h3e5c94fe,
32'hbe91858f,
32'hbc91ddce,
32'hbe4da906,
32'hbd32232e,
32'hbe0b79ca,
32'h3ebe50a7,
32'h3ece3149,
32'hbfa83574,
32'h3d41aa86,
32'h3f0ada50,
32'hbdf2a474,
32'h3ea85ae7,
32'h3f0b5df7,
32'h3e3b0837,
32'h3eac89a0,
32'hbe117956,
32'hbd50ffe0,
32'h3d3630dc,
32'h3f28df0a,
32'h3ddf4c41,
32'h3ce18a34,
32'h3f2322d0,
32'h3eda7482,
32'hbe5d4afa,
32'hbe709701,
32'hbdbfce75,
32'hbf37cc16,
32'h3e5389ce,
32'h3eec2f87,
32'h3f169734,
32'hbf081ae3,
32'hbe472bcd,
32'hbd51615d,
32'hbc2627a1,
32'hbceb602b,
32'h3ea8e5e5,
32'h3f05a356,
32'hbdca9811,
32'h3e9eb801,
32'h3d3a938c,
32'h3e6b6b2f,
32'h3e947f24,
32'h3f282691,
32'h3e849a37,
32'h3d81b4f7,
32'hbe70a328,
32'hbcdb6c75,
32'h3ceccbaa,
32'h3ee3a02a,
32'h3df9fa9f,
32'h3dfff821,
32'h3f284d2c,
32'h3ef1daf4,
32'hbe38fccf,
32'h3b752188,
32'hbe64f076,
32'hbdb6fe63,
32'h3ea07f37,
32'h3f2ff8e7,
32'h3f355593,
32'hbe8d574f,
32'hbe4526fc,
32'hbcbd92e1,
32'hbc8fdabd,
32'hbe502214,
32'h3e5c6f55,
32'h3eafda6e,
32'h3e79a861,
32'h3edbfbc5,
32'hbe6d5182,
32'h3ec98c94,
32'hbb162bc3,
32'h3edf7316,
32'h3efcaaa9,
32'hbe8b08c2,
32'h3d7bc089,
32'hbb270aa1,
32'hbd5f1ebe,
32'h3ea428fc,
32'hbdc7ea6a,
32'h3e3387c8,
32'h3f05bbfa,
32'h3e9b58cc,
32'hbed4f2cf,
32'h3e1d997e,
32'hbea8f5d0,
32'hbeecb149,
32'h3ecdde09,
32'h3f40abe8,
32'h3f28dc63,
32'hbedbec6c,
32'hbddd6a58,
32'h3e538660,
32'h3eb20d1f,
32'hbeb3856d,
32'h3e53fe43,
32'h3e1eaf49,
32'h3e498f3f,
32'h3f031972,
32'hbe603e03,
32'hbd47cfc5,
32'h3e0a7ab1,
32'h3df0fb8b,
32'h3e5a1722,
32'hbe517a64,
32'h3eb69479,
32'hbe11d028,
32'hbcd0c47a,
32'h3ea54704,
32'hbbd5c2ca,
32'h3eb66892,
32'h3eb4bc1a,
32'h3dacc635,
32'hbdea2c06,
32'hbe29d552,
32'h3d814c5d,
32'hbe9b7bdb,
32'h3e8491ed,
32'hbcdf6b07,
32'h3e8efe14,
32'hbe212b2c,
32'hbdee1669,
32'h3e042bc8,
32'h3eda093c,
32'hbe9a0303,
32'h3e662ced,
32'hbef6b939,
32'h3eec03c9,
32'h3e883477,
32'hbb157ba0,
32'hbee605b4,
32'h3eb07353,
32'h3dbc86f4,
32'hbd397ca8,
32'h3d792fab,
32'h3ee8d934,
32'hbd487c0d,
32'h3b9bab73,
32'h3ef42619,
32'h3da4dfc6,
32'h3e77221d,
32'h3d227e89,
32'hbeb92348,
32'hbd0ed0d5,
32'h3e87d355,
32'h3e4e6855,
32'hbd4225a4,
32'hbdb59d88,
32'h3cecc13b,
32'h3e6a1cd9,
32'h3e02b9c3,
32'h3e25489b,
32'hbec4603f,
32'hbdba3af6,
32'hbf0bf3ca,
32'h3dedd754,
32'hbee68533,
32'hbdee311c,
32'hbccafd1d,
32'hbe02e305,
32'hbe95b826,
32'h3e03a9c4,
32'hbe08cbdf,
32'h3d9249d4,
32'hbdeffa18,
32'h3dd7b07b,
32'hbd9659de,
32'hbc254325,
32'h3e1eb4c4,
32'h3eab614b,
32'h3d4ff524,
32'hbd8aef10,
32'hbf2e9065,
32'hbd7d2c37,
32'h3e5f382f,
32'h3e62d078,
32'hbe1e5530,
32'h3dc8ea24,
32'h3eb838db,
32'h3c949e91,
32'hbd1f343c,
32'hbe16e2ab,
32'hbd25e350,
32'h3e9d5f27,
32'hbe74f90d,
32'h3e89522c,
32'hbf1f3248,
32'hbdb9d1fc,
32'hbde62ef5,
32'hbd98753c,
32'hbe535d91,
32'h3e165cf8,
32'hbdf3a249,
32'h3cbb8bde,
32'h3e0d05e8,
32'hbae8dcc3,
32'hbd26d2cf,
32'h3cd0c6a5,
32'h3e143fb0,
32'h3e476ebe,
32'hbe025466,
32'hbdf58193,
32'hbcf83d56,
32'hbcec4d67,
32'hbdccad45,
32'h3e7fc1ef,
32'hbe95f933,
32'h3e29ebf7,
32'h3e3c28ca,
32'h3e0465b6,
32'h3d308b81,
32'hbedcd574,
32'h3d9546ec,
32'h3ed19136,
32'hbdff96fd,
32'h3bcdf660,
32'h3eb31c82,
32'h3d68fa81,
32'hbe13319d,
32'h3dada0c5,
32'hbe415e77,
32'hbdf251ac,
32'h3e1d8cf2,
32'h3d8e1db0,
32'h3e39b93a,
32'hbda6ce63,
32'hbd430791,
32'h3d93b7d4,
32'h3e006df2,
32'hbb5bd790,
32'hbd28dff9,
32'hbe015b7d,
32'h3e7cfcd4,
32'hbe07be08,
32'h3c1018e0,
32'hbd3c6c23,
32'hbeb7a238,
32'h3e238ab7,
32'h3dc3966f,
32'h3e989a86,
32'h3e066a53,
32'hbe6225ca,
32'h3e325199,
32'h3e600b06,
32'h3e259a96,
32'hbd409772,
32'hbf8125bc,
32'h3e2c7581,
32'h3dd03387,
32'hbda0330c,
32'hbf430d84,
32'h3d96bf63,
32'h3e9e4725,
32'hbe4dca00,
32'h3c54a14e,
32'h3e644e0f,
32'h3c89357e,
32'hbd7f9f13,
32'hbdeb27f1,
32'h3e65b76d,
32'h3e18d837,
32'hbe95d20a,
32'h3f1c4b8f,
32'hbdeb5235,
32'hbee13022,
32'h3e4ef100,
32'hbf0c897d,
32'h3da9b2cf,
32'h3ebc12f9,
32'h3e6f509f,
32'h3e02b7f4,
32'hbf2d8124,
32'h3e989cda,
32'h3e929385,
32'h3deacb82,
32'hbe4bc42a,
32'h3e88f55f,
32'h3d1fafd3,
32'h3e78d581,
32'hbdf14245,
32'hbec40314,
32'hbe3efc73,
32'h3ec30fd2,
32'hbec3f5a5,
32'h3dd39abb,
32'h3e2b41ad,
32'h3d27f67e,
32'h3d168278,
32'h3df26668,
32'h3d3f60b4,
32'h3d21c9f6,
32'hbe1a44c7,
32'h3df5ca6a,
32'hbbbe6a71,
32'h3e42fab2,
32'hbc8129f1,
32'hbf590ca7,
32'h3c54c27c,
32'hbe56397e,
32'h3e3ab4b4,
32'h3d5be415,
32'h3e741d1b,
32'h3eb1cd5d,
32'h3d87e16f,
32'hbd1c8ce6,
32'h3d659334,
32'hbee682bd,
32'h3db0872c,
32'h3cc0fd8a,
32'h3d7e5e62,
32'hbdd4d52f,
32'h3e033fe7,
32'h3e38d383,
32'hbeca7f34,
32'hbd405125,
32'hbe8316cd,
32'hbde7389c,
32'hbd1ddf6e,
32'h3e9422e1,
32'h3d8e5793,
32'hbe3a02b3,
32'hbe6c2c3c,
32'h3e923f1f,
32'hbd75e24f,
32'hbe8a9e56,
32'hbe8fd46b,
32'hbf4e201d,
32'h3c8106f2,
32'hbe283101,
32'h3e5e39d7,
32'h3dc420a2,
32'hbe6b73cb,
32'h3d69549e,
32'h3dd21ea9,
32'hbb304584,
32'hbe03c9a5,
32'h3bd15f67,
32'hbeee12a1,
32'hbdfe6260,
32'h3e8d745e,
32'h3ddd058b,
32'h3dff35de,
32'h3eba48e3,
32'hbf5e3467,
32'h3ef51eec,
32'h3ec5183f,
32'hbb943b7f,
32'hbcec6025,
32'h3d53b7a8,
32'h3e1b6186,
32'h3d1fa245,
32'hbe5ae227,
32'h3efbd427,
32'hb8a32e8f,
32'hbebb039c,
32'h3cd6f2ca,
32'hbf895aa6,
32'h3dd1dca8,
32'hbe4e5f4b,
32'h3e57dcf6,
32'h3e9ee733,
32'hbf55d079,
32'h3da11eb7,
32'hbec92676,
32'h3d8baf9e,
32'h3e1a6ea7,
32'hbee6374b,
32'hbe882834,
32'hbe4ab367,
32'h3f140485,
32'h3e002487,
32'h3eb90976,
32'h3eaf4d85,
32'hbf4116f5,
32'h3f5dce3f,
32'hbdb91588,
32'h3d24c425,
32'hbba281af,
32'h3d4f855d,
32'h3c9e24f3,
32'hbe8b17fe,
32'hbdba72bb,
32'h3eaad077,
32'h3e9e24ed,
32'hbf05f4bb,
32'hbf1fc156,
32'hc00f77bc,
32'hbc131e1c,
32'h3e886127,
32'h3e391367,
32'h3e6d728c,
32'hbf7f2d60,
32'h3e7e92db,
32'hbe2c970a,
32'h3d503b20,
32'hbf17c292,
32'hbee5eb24,
32'hbf8bd742,
32'hbeaa44db,
32'hbe09955b,
32'hbec573e8,
32'h3eb6aadd,
32'h3ec4ebce,
32'h3d67e8ba,
32'h3f028a3a,
32'h3e28c4ce,
32'hbdffd904,
32'hbd4e5138,
32'hbe811d17,
32'hbe824490,
32'hbdf356c8,
32'hbdbed1c7,
32'h3d5c665b,
32'h3e451ebf,
32'hbf14053c,
32'h3dc17fab,
32'hbf9fff21,
32'h3dae4b86,
32'h3e8ea085,
32'hbe0ef677,
32'h3c2696cb,
32'hbd871a2d,
32'h3e531f8f,
32'h3eade4e1,
32'h3e960678,
32'hbe7f738d,
32'hbc9fb801,
32'hbf949ee4,
32'hbf05ad69,
32'hbdf963b5,
32'hbf3461e6,
32'h3f9db2f2,
32'h3cbc9d78,
32'h3ed7eb78,
32'h3e02414a,
32'hbede3aa9,
32'h3d1bf955,
32'hbc77bda4,
32'hbe8960f0,
32'hbeacb089,
32'h3e9deb2b,
32'hbd95b358,
32'h3f35f85c,
32'h3ea7919d,
32'hbf4ab1d1,
32'hbe8b39b7,
32'hbf57b6d3,
32'h3de3750f,
32'hbfbfc19c,
32'hbcb597bd,
32'hbf1b174c,
32'h3e23b946,
32'h3de6f664,
32'hbf12012b,
32'h3eea69cb,
32'hbdcb78f4,
32'h3f629055,
32'hbe4edc14,
32'h3f52ff5a,
32'hbf3d9791,
32'hbc19a1df,
32'h3f64a9bb,
32'h3c749d8b,
32'hba4f7b9c,
32'h3de7a758,
32'hbec1dda3,
32'hbc439b06,
32'h3ce6d279,
32'h3b127e97,
32'hbe266a2f,
32'h3f549914,
32'hbade9203,
32'h3f053ab2,
32'hbf83eca3,
32'h3e6e12f2,
32'hbf3fa65e,
32'hbf516bb4,
32'hbec44ea8,
32'hbe2abac3,
32'h3db37361,
32'hbe93d754,
32'h3e04f54f,
32'h3de09763,
32'hbf2617e2,
32'h3e34365d,
32'hbe60adbe,
32'h3f15f172,
32'h3d0ba7b1,
32'h3fc2c168,
32'hbf3313bc,
32'h3b57ae77,
32'h3c532d1b,
32'h3f1ca9db,
32'h3e7849f6,
32'h3f5dc516,
32'h3e727e6d,
32'hbd1d65eb,
32'h3d9b4e3a,
32'hbece86a5,
32'h3ee0d73b,
32'h3e8ba04a,
32'h3d9c0476,
32'h3fc638db,
32'h3d08292d,
32'h3d0a32fe,
32'hbe9435d4,
32'h3efa7605,
32'hbf20b044,
32'hbeb0b27b,
32'hbf6e6f9e,
32'h3f70b74f,
32'h3e897c56,
32'h3f7ba778,
32'h3e7e04c4,
32'h3f95d0e8,
32'hbf2072be,
32'h3c0fc770,
32'hbd40ed34,
32'hbda967ad,
32'hbe682201,
32'hbcca0ca3,
32'hbe24e1da,
32'h3f3f6507,
32'h3d6de811,
32'h3d80d47e,
32'h3e015e06,
32'h3beec549,
32'hbccbe129,
32'hbe395c6c,
32'h3f41ef62,
32'h3c019f81,
32'hbe860070,
32'h3f4b95c4,
32'h3dae881a,
32'h3c74f9ab,
32'h3b826a00,
32'h3e12a1e0,
32'hbecf8d4a,
32'hbe52301f,
32'hbf3bb8ec,
32'h3ee96f45,
32'hbdb04e55,
32'h3f52cc93,
32'hbd63ea55,
32'h3d33033e,
32'hbed99ced,
32'hbd87e554,
32'hbd02af8f,
32'hbdaebfd5,
32'hbd344c7c,
32'hbdab85f3,
32'hbd8b0697,
32'h3d85f9bd,
32'hbbc27591,
32'h3d5f8068,
32'h3cc87871,
32'hbc6c74eb,
32'h3d948533,
32'hbcf4c137,
32'hbd9eb3c1,
32'hbc822590,
32'hbd643753,
32'hbcab4a4a,
32'h3d82634c,
32'h3b142039,
32'hbc8e85d8,
32'h3d9bf6bd,
32'h3d3bfe0c,
32'h3d07448a,
32'hbd90f4aa,
32'h3d4bd53f,
32'h3c801deb,
32'h3d40e373,
32'h3daac2d5,
32'hbc33ceea,
32'h3bd6b14b,
32'hbcaeaf8b,
32'hbc0685dc,
32'h3e56c109,
32'h3d7a96cf,
32'hbd366253,
32'hbe9daad9,
32'h3e5f9cba,
32'hbdc32266,
32'hbba01f6e,
32'h3da35a5c,
32'hbcdcf4f3,
32'hbd1649c6,
32'hbec19932,
32'h3e8b07f6,
32'h3e9123d2,
32'h3dabe559,
32'hbcb7f196,
32'h3d045a03,
32'h3e9cd33c,
32'h3ce427a8,
32'h3e183d3c,
32'h3ee8ba4a,
32'h3d26db48,
32'hbd89cc49,
32'h3dc49231,
32'h3d341ac1,
32'hbcde5acf,
32'h3d5783c3,
32'h3d32688b,
32'hbe16a6ee,
32'h3e181064,
32'h3f5ab59c,
32'h3e31d0ff,
32'h3f6301ab,
32'hbeccf29c,
32'h3fbf5cc4,
32'hbe51dc7b,
32'hbda85d75,
32'hbe15b782,
32'hbec7a426,
32'h3d490343,
32'h3ca392a7,
32'hbeddf3f7,
32'h3efa8269,
32'hbdcf1115,
32'h3e2b54aa,
32'hbdbdbefa,
32'h3f125872,
32'h3e31ade3,
32'h3e24048f,
32'hbf133809,
32'h3f0230b7,
32'h3cdf74ca,
32'hbe07fb06,
32'hbf1f9ab5,
32'h3f69aa2b,
32'hbd9ead04,
32'h3c42cb41,
32'hbdaf08d4,
32'h3e3c563d,
32'hbe296027,
32'hbf5576dc,
32'h3da1ce18,
32'hbd815c43,
32'hbeb3504a,
32'h3c653c8c,
32'h3d687dd5,
32'h3f291946,
32'h3eacb38e,
32'hbec14044,
32'hbcab6bac,
32'h3ce97bf5,
32'h3dbe052c,
32'h3e106210,
32'h3d29a78d,
32'h3d0c7c1c,
32'h3de8ea36,
32'h3d01ec67,
32'hbe06d295,
32'h3f0a73cb,
32'hbe5f31a0,
32'h3e305b9a,
32'hbebf534b,
32'hbe86788e,
32'h3f6f5246,
32'h3ccf7f9b,
32'h3efa0c20,
32'hbe07da34,
32'hbd19f956,
32'h3e6d59ad,
32'h3f180251,
32'hbf1ce9cb,
32'hbcf01949,
32'hbcdd445d,
32'hbf5b896f,
32'hbdd4f8ab,
32'h3d1cee71,
32'h3d3a9094,
32'h3e40a23c,
32'hbf23d0e1,
32'hbd670b4b,
32'hbd0604e3,
32'h3f00ea48,
32'h3aff98ce,
32'hbd456b1c,
32'hbe116f08,
32'hbcd4aced,
32'hbf6af198,
32'hbfccd2aa,
32'h3cebc83f,
32'h3ea58fa2,
32'hbe24c28e,
32'hbf6dc9e9,
32'hb933609c,
32'h3e95749c,
32'hbeaf3991,
32'hbb91b35c,
32'h3edce705,
32'hbd504d81,
32'hbe4e5b8a,
32'hbea97ca7,
32'hbeaa62c9,
32'h3ead45df,
32'h3dcc8dda,
32'hbf0044bb,
32'h3e20e535,
32'h3e24baa6,
32'hbe1ef22d,
32'h3def1626,
32'hbfae874f,
32'h39ec31d3,
32'hbd3e9efd,
32'h3e307a77,
32'h3eb1e951,
32'h3e357612,
32'hbe497973,
32'h3eaba404,
32'hbea9cdd1,
32'hbef5458a,
32'hbd44553a,
32'h3df65709,
32'hbe4abc41,
32'hbf2bde69,
32'h3d894271,
32'h3eef0706,
32'hbf0a4beb,
32'h3da17361,
32'h3e6dfdc6,
32'h3ef22c0e,
32'hbf37f4d3,
32'hbc394051,
32'hbf2ae80b,
32'h3e3d6011,
32'hbb963f34,
32'hbf1f00c8,
32'hbe3e1d19,
32'h3c580b11,
32'hbddf046e,
32'hbd528c44,
32'hbf487014,
32'hbd11eac6,
32'hbc805210,
32'hbe5802e8,
32'h3cf85388,
32'h3ddcd6a5,
32'hbc6032f8,
32'hbead7f9c,
32'hbec6fdf8,
32'hbeab5342,
32'h3e00a89d,
32'hbffef3d1,
32'h3e9f32e6,
32'h3e33c060,
32'hbd67e705,
32'h3df3f492,
32'h3f18d326,
32'h3e7a5b74,
32'h3ee84985,
32'hbed06139,
32'h3c0c86ed,
32'h3e01772e,
32'hbf63d5b1,
32'h3dbb66cf,
32'h3df0beac,
32'hbe3d0451,
32'hbe17bd46,
32'h3dbb4ca2,
32'hbde3324d,
32'hbddd59f6,
32'hbf211eb9,
32'h3c61791c,
32'hbdca677a,
32'h3bcc01e6,
32'h3e898090,
32'h3e25d305,
32'h3d0bd2a8,
32'h3e73fc18,
32'hbeaba944,
32'hbf25dd5e,
32'h3e3a6562,
32'hbfbcd198,
32'h3dbf60e7,
32'hbc763771,
32'h3c512f4a,
32'hbdbbd25c,
32'h3f402aee,
32'h3e9d4e75,
32'h3e617f57,
32'hbe2165ce,
32'hbd85b66a,
32'h3e081e9c,
32'hbf755486,
32'h3ea72088,
32'hbc420e2c,
32'h3e3f66df,
32'h3dddf813,
32'h3c5c1102,
32'hb900f06a,
32'hbe73a59c,
32'hbef47b1a,
32'h3c6f71c0,
32'h3d1d5fc5,
32'h3c1845af,
32'h3ebb8a48,
32'h3f054e2b,
32'hbd214004,
32'h3d78751f,
32'hbef97895,
32'hbf8ee36f,
32'hbb3ad189,
32'hbe9fb5ec,
32'h3dd44b74,
32'h3d034586,
32'h3e397e23,
32'h3defc36e,
32'hbc0ad7e5,
32'h3e8e4f5b,
32'h3e383371,
32'hbe37acdc,
32'hbe51ecf2,
32'h3e18dc7f,
32'hbfba92f2,
32'hbdd41715,
32'h3f0387da,
32'h3c4bae5b,
32'h3e9d22b6,
32'h3d9c1c38,
32'hbbe05430,
32'hbe6e3de4,
32'h3ee65b8c,
32'hbe0ccfe8,
32'hbdecfbb7,
32'h3cea9fdb,
32'h3e931f42,
32'h3dfbf2ff,
32'hbd9a0bc4,
32'h3db8dd36,
32'hbf5039e9,
32'hbf447f28,
32'hbf19788f,
32'h3f1d4097,
32'h3cfe325a,
32'hbe2251ec,
32'h3e5eda05,
32'h3dc7f088,
32'hbe883f1a,
32'h3e428f37,
32'hbd4ea7dd,
32'hbe1c1320,
32'h3d9cd556,
32'h3e1d5a06,
32'hbcb775fb,
32'h3dab2bc5,
32'h3ee8c993,
32'h3d686c9d,
32'h3ec708b2,
32'h3d2399a3,
32'h3d3685ba,
32'h3e44b18e,
32'hbe65ede0,
32'hbdd689a3,
32'hbd02721a,
32'h3edefd6c,
32'h3df7b3c4,
32'h3ddac089,
32'h3c4a1f49,
32'h3e23f2ae,
32'hbe69488a,
32'hbf812a0d,
32'hbed1875f,
32'hbb96160d,
32'h3dc13e9d,
32'hbc245669,
32'h3e8580d5,
32'hbdeec2ab,
32'hbe7d1f39,
32'h3e4177f8,
32'h3e09e09e,
32'h3e1fac33,
32'h3eb0b59d,
32'h3ed96372,
32'h3cb94831,
32'h3ed85a48,
32'h3ed5334c,
32'h3e8e84ec,
32'h3e5df073,
32'hbd473bdb,
32'h3dd02c7e,
32'h3e1d788c,
32'h3c8b726c,
32'hbdcedc58,
32'h3d392fe1,
32'h3eea69e4,
32'h3e311ca3,
32'h3dd90fb8,
32'hbd12cd5f,
32'h3da7810d,
32'hbe9691f8,
32'hbee54af2,
32'hbeaffc27,
32'h3adadb25,
32'h3e9c883f,
32'h3ea424b8,
32'h3e95f6a8,
32'hbe96f8b5,
32'hbd15886c,
32'h3e7a474c,
32'h3e3e6d25,
32'h3dfd1a99,
32'h3de6034d,
32'h3e963027,
32'hbe71b533,
32'h3ea5ad33,
32'h3e4c9cbc,
32'h3e12ea35,
32'h3cbe5ca9,
32'h3cec1b86,
32'hbce2abf1,
32'h3dec5d78,
32'h3ee3fc2d,
32'hbd586b56,
32'h3c5006e5,
32'h3eb1d2dc,
32'hbddf5243,
32'h3e0585e5,
32'h3c201928,
32'h3d626e13,
32'hbd858093,
32'hbe6b1bf8,
32'hbe3fab21,
32'h3dd4d461,
32'h3dc94bd7,
32'h3e5f2174,
32'h3ebf1818,
32'hbe269a94,
32'h3c907508,
32'h3d2d4435,
32'h3de8f132,
32'hbeb95656,
32'h3ebdf087,
32'hbe90466e,
32'h3e867418,
32'h3e19fdea,
32'h3d7ed3c2,
32'hbd90f55e,
32'hbd71bfa2,
32'h3e34c8dc,
32'h3ea80a77,
32'hbe91c2ea,
32'h3e28a5e2,
32'hbd9033bd,
32'hbd71c6be,
32'h3e4922cf,
32'hbec5e3e3,
32'h3d73bf5c,
32'h3dbf63d7,
32'h3d235ff6,
32'h3e3adb75,
32'hbe5819c6,
32'hbe056e8b,
32'h3d4f4e06,
32'h3e985bc8,
32'h3f14c444,
32'h3e2c8903,
32'hbe506c67,
32'hbea2d717,
32'hbd0c3142,
32'h3bc67043,
32'hbed8ce58,
32'h3ee55c43,
32'hbedf2544,
32'h3eca7ad3,
32'h3ceffc38,
32'hbe30f161,
32'hbf038559,
32'h3de6cd6e,
32'h3d4b7160,
32'h3d9a270e,
32'hbe8315a3,
32'h3e325eae,
32'hbcced8fe,
32'h3d7cb1a2,
32'h3e9fc2a5,
32'hbe0d6f0f,
32'h3e543df6,
32'hbe41499a,
32'hbda9131b,
32'hbdbfc510,
32'hbd499e4f,
32'h3b8c7044,
32'h3e6dd78c,
32'h3d4cfbe0,
32'h3ea08901,
32'hbe1b77a3,
32'hbd7f1721,
32'h3e88e747,
32'h3ccfdf4a,
32'hbe0e9e6d,
32'hbf5f6dc9,
32'h3edcb7d5,
32'hbf14c7bc,
32'hbda8e84d,
32'hbca87a8e,
32'hbdf496ff,
32'hbf2097ba,
32'hbd5161c6,
32'hbdb88d32,
32'h3dc9206b,
32'hbed56ec1,
32'h3cef0b04,
32'hbcfffe5f,
32'hbd5c9b75,
32'hbd2fcb03,
32'hbd056bde,
32'h3e2f55e0,
32'hbdab02c6,
32'h3e93797e,
32'h3c644156,
32'hbec97c4e,
32'h3e6149d5,
32'hbe7df3bf,
32'h3e5a41d0,
32'h3ec90c43,
32'h3c9967ab,
32'hbdaeaad4,
32'h3d484178,
32'h3eb4cbdc,
32'hbd53507c,
32'hbf3f055b,
32'h3e708d73,
32'hbf1a4ed7,
32'h3cc2249b,
32'h3d03572a,
32'hbdad1572,
32'hbf199be7,
32'h3d9c90d8,
32'hbe103b38,
32'h3c10191d,
32'hbeb12f3f,
32'h3ea348bc,
32'hbc5c172f,
32'hbb6c2372,
32'hbdd06149,
32'h3e71eee8,
32'h3e83ebbb,
32'h3daaf4ef,
32'h3e58b5a7,
32'hbacb52bb,
32'h3d23e9d1,
32'hbd1550f6,
32'hbd469021,
32'h3e2c268f,
32'h3c93b9fe,
32'hbd0945a2,
32'hbdb63eb8,
32'hbe9bad76,
32'h3e444ceb,
32'h3e60b1a0,
32'hbedc2162,
32'h3d88e59f,
32'hbda93533,
32'hbd909ce3,
32'hbced6d9c,
32'h3e444be8,
32'hbf72a92e,
32'h3e9a84fe,
32'hbe652569,
32'hbe9dd1c1,
32'hbf0b4875,
32'h3e0b45bc,
32'hbd582b38,
32'hbde16cf6,
32'hbc044e3b,
32'hbd8b80f9,
32'hbe024d75,
32'h3d834b7e,
32'h3e8c1833,
32'h3c354abd,
32'hbeed227a,
32'h3de29c72,
32'hbeb8db94,
32'h3dcd97f1,
32'h3d803948,
32'hbe327354,
32'hbe6b3d8e,
32'hbe9192c9,
32'h3e42dba9,
32'hbe60fe74,
32'hbe233ec7,
32'hbd74cafc,
32'hbf2f34c2,
32'hbd344084,
32'hbd4df1be,
32'hbd7e5949,
32'hbf19a93b,
32'h3e46edf0,
32'h3d8c7f15,
32'hbe72f86c,
32'hbeb8c2c6,
32'h3eadc5ac,
32'hbd04dfdf,
32'hbd78472e,
32'h3d0c5b9e,
32'h3dd39e57,
32'hbe6b7b42,
32'hbc5ef042,
32'h3d23df4d,
32'h3d76d6e8,
32'hbed5b7f9,
32'h3ee97a75,
32'hbe5d9b39,
32'hbc3ca450,
32'h3e5268e3,
32'hbe6f7e84,
32'h3e830a78,
32'hbf9b6e49,
32'h3dceb350,
32'hbd414bd8,
32'hbe986b64,
32'h3d94132d,
32'hbeb22d39,
32'hbe65cc87,
32'h3cc90649,
32'hbe776f49,
32'hbcb8495d,
32'hbe27ca8d,
32'hbe04668b,
32'hbecbdeb9,
32'hbeb2d78e,
32'h3db07992,
32'h3ca648d9,
32'hbd2c29bc,
32'hbdb1aec1,
32'h3dfbecd5,
32'hbccef55a,
32'hbdbf8498,
32'hbc39c961,
32'h3e3652f6,
32'hbec57755,
32'h3e689388,
32'hbf0c3748,
32'hbe2e9e22,
32'h3e5c13c4,
32'hbe2b158e,
32'hbe0fa462,
32'hbf35c7c2,
32'h3e5c7d8a,
32'h3e1f727b,
32'hbe59ab7b,
32'h3e2288b4,
32'hbffce1e1,
32'hbf07efb7,
32'h3e34ddbb,
32'hbed37a52,
32'h3de98a9f,
32'hbe539348,
32'hbd224661,
32'hbeec21ef,
32'h3e3b6a3a,
32'hbe095d93,
32'h3c42acf3,
32'hbdb8d7b7,
32'hbdb76da1,
32'h3d1b11fa,
32'h3eb6c696,
32'h3b656ccc,
32'hbdfb61ed,
32'h3e26336d,
32'hbf469ea0,
32'h3ceb3d5d,
32'hbf935f70,
32'h3e20bb67,
32'hbc9fd83a,
32'h3a949c84,
32'h3d624b5d,
32'hbfbfb866,
32'h3eedb7c5,
32'h3ce9762f,
32'hbe3430f6,
32'h3da7e581,
32'hbf3a5fc8,
32'hbf536b6c,
32'hbd43b4ec,
32'h3bb9eadc,
32'h3e193711,
32'h3ea9b1d0,
32'h3e722c98,
32'hbf4f306c,
32'h3e2f98e1,
32'hbca84e1b,
32'h3d3a4906,
32'hbd10d230,
32'hbdcd8a1d,
32'hbeda3493,
32'h3debc6fe,
32'h3e061dfa,
32'hbd7d94b1,
32'hbe0b004c,
32'hbf23712a,
32'h3e30d41c,
32'hbf6fad43,
32'h3e6ff12f,
32'hbe51eff5,
32'h3e5c3332,
32'hbd56679b,
32'hbf974824,
32'h3ed55aec,
32'h3cc041d4,
32'hbe93e085,
32'hbe0dcbb6,
32'hbf05829a,
32'hbe14be1e,
32'h3e09660b,
32'hbdd9c29b,
32'h3e4d1c5e,
32'hbd7d51bc,
32'h3ecf0e3b,
32'hbf054815,
32'h3e8e8c13,
32'hbe992071,
32'hbc290f8d,
32'hbd07e6bf,
32'hbe8a7c56,
32'hbeb37e20,
32'hbda88568,
32'h3e4e0b0e,
32'h3eaf3658,
32'h3d8b19b7,
32'hbebc58f4,
32'h3dee7059,
32'hbf93fc90,
32'hbc8b6588,
32'h3d8b5ebd,
32'h3e7edcd2,
32'hbf181b6a,
32'hbecf9f5b,
32'h3e9c2209,
32'h3d8ded52,
32'h3dccf2da,
32'hbf365f02,
32'h3e71c2e2,
32'hbee573ac,
32'hbc968974,
32'hbde12daa,
32'h3ddf5547,
32'h3d9376d7,
32'hbeb03b93,
32'hbdcb13b3,
32'h3ecc4311,
32'h3e20df7e,
32'hbdd733ac,
32'hbb260546,
32'hbefc8594,
32'h3d1b7c75,
32'h3ed0e663,
32'h3e3b34d0,
32'h3e382202,
32'h3dea9e5f,
32'hbf7e07dc,
32'h3f2fa926,
32'hbe1b9c9c,
32'h3e85847a,
32'h3f804490,
32'hbe7f6012,
32'hbf1427a7,
32'hbf0cd238,
32'h3e876e78,
32'h3f4174b0,
32'hbe662b65,
32'hbf4983f8,
32'h3f1635f2,
32'hbeab0aa3,
32'hbebab638,
32'hbd5cd8d5,
32'hbea5bd54,
32'h3fc211d5,
32'h3d35f6d1,
32'hbbacdc62,
32'h3e8a11fb,
32'h3de272ff,
32'h3cec1539,
32'h3b4e0889,
32'hbe9843fa,
32'h3f166081,
32'h3f2bc4df,
32'hbf0c19a0,
32'h3edc00d1,
32'hbe3e5b46,
32'hbda239a4,
32'h3f013a73,
32'hbee1ba1b,
32'hbe3c83c1,
32'hbfa75502,
32'hbf042bfc,
32'hbebb6314,
32'hba9b5bef,
32'hbdad8faa,
32'hbeb9049b,
32'h3f49d39b,
32'hbf0f84c0,
32'h3f84ff6d,
32'hbe0ca2ba,
32'h3f9b868f,
32'hbe580374,
32'hbe9acc32,
32'hbf0c4102,
32'h3f1e6b09,
32'hbd2bf2b4,
32'hbe4233ae,
32'hbeab9623,
32'hbaa97c09,
32'hbca0119b,
32'hbe821bfb,
32'h3e85cff1,
32'h3f3c1a39,
32'hbe3e684c,
32'h3efad5fa,
32'hbeafc164,
32'h3f4005f5,
32'h3c641655,
32'hbe6e3349,
32'h3e316995,
32'hbf83dc03,
32'h3ea1a76d,
32'hbee9d4ea,
32'hbd9d4752,
32'h3efa3bd7,
32'hbecec9f8,
32'h3f0bd5cc,
32'hbe0b3d83,
32'h3f23eb19,
32'h3cd212ef,
32'h3fe93e4f,
32'h3f17b657,
32'hbdf1e91f,
32'h3e1e137f,
32'h3f1963d5,
32'hbd5decf0,
32'h3ffc2a98,
32'hbc6eb2e1,
32'hbdbf4a25,
32'h3d73df8a,
32'h3f02a5fa,
32'h3fb79d18,
32'h3ebb6625,
32'hbeaf0720,
32'h3f908e0e,
32'h3da6f729,
32'hbf3549bc,
32'hbf303589,
32'hbe6a49f1,
32'hbeae71ec,
32'hbf2b8490,
32'hbf60997d,
32'h3fa047fa,
32'h3e81f01e,
32'h3ec41ad8,
32'hbd3e1503,
32'h3f3f10d7,
32'hbf15a68d,
32'h3c4e583e,
32'hbcf78f28,
32'h3cc1afea,
32'h3cc279f9,
32'h3b83a893,
32'hbb35962d,
32'h3c8a3574,
32'h3c80eb27,
32'h3d4748cd,
32'h3bf358f5,
32'hbd1ff37a,
32'h3de81232,
32'hbd0ef8b2,
32'h3d441980,
32'h3c9f9928,
32'h3bd4cc06,
32'hbbc70186,
32'hba30f816,
32'hbd2f0ecf,
32'h3cfbf157,
32'hbe0f1c8c,
32'h3e653379,
32'hbd76937e,
32'hbd2b26f7,
32'hbc8b60aa,
32'h3cf9b14c,
32'h3ea8c7f7,
32'h3e09f25a,
32'hbc0a7ab0,
32'h3dc9c0cd,
32'hbd566b38,
32'h3d64a6eb,
32'hbd84f513,
32'hbd8d6926,
32'hbd94f99c,
32'hbd58f63c,
32'h3c46d609,
32'h3dbf9260,
32'h3caaf0e6,
32'h3d818f17,
32'hbd9a2ade,
32'hbd5a3c60,
32'h3d8898ae,
32'h3cbdd0a2,
32'h3d1148c4,
32'h3df2b5c3,
32'hbb4524df,
32'hbd0a3050,
32'hbd012fc5,
32'hbce30373,
32'hbd477d8d,
32'h3d81a230,
32'hbd174790,
32'hbb62783a,
32'hbabfd0d9,
32'h3c4b6c2d,
32'h3e0f6442,
32'hbd8ef445,
32'h3d61dafe,
32'h3d2d4754,
32'hbdd5b664,
32'h3d89e7d0,
32'h3e22c1a7,
32'hbdcfdba9,
32'h3cbc8ed8,
32'hbe82dc33,
32'h3e926752,
32'h3e41f0d9,
32'h3d3783c8,
32'h3d4c5767,
32'h3c1a3245,
32'hbabe5c00,
32'hbeb8bcf7,
32'h3e8a198c,
32'h3eb6fd07,
32'h3ecd2b6e,
32'hbccaea1b,
32'h3d0f5979,
32'h3d68d97f,
32'h3b888098,
32'h3e146ffb,
32'h3f0db231,
32'h3d43d805,
32'hbe233e58,
32'h3ec920e3,
32'hbc2a105f,
32'h3e30c942,
32'h3cf95158,
32'hbd8665eb,
32'h3d4da654,
32'hbe214378,
32'h3e326bc1,
32'h3e5c740c,
32'hbe959b4d,
32'hbd3d7b4e,
32'hbf17730d,
32'h3e1925b0,
32'h3e364589,
32'h3f011a84,
32'hbdc8e08e,
32'hbcc8b366,
32'hbd131355,
32'hbf4487d5,
32'h3f5f38b6,
32'h3d971be3,
32'h3dbe0559,
32'h3ededd50,
32'h3ef68f10,
32'h3d64072e,
32'h3df012d3,
32'h3daefce6,
32'h3f42516b,
32'h3dc314a0,
32'h3d25002f,
32'hbdd3f582,
32'h3c39442f,
32'hbf220f9e,
32'h3e74c643,
32'hbdc38e53,
32'hbdcf4625,
32'hbd707e97,
32'hbf94ae98,
32'hbf812d49,
32'hbf223316,
32'h3f03c2be,
32'hbe931280,
32'hbd54bd09,
32'h3d79ffac,
32'h3f293ffe,
32'h3d4c9f80,
32'hbca1529d,
32'h3c0db46c,
32'h3e4203bf,
32'h3f341078,
32'h3db374e9,
32'hbee9e83b,
32'h3f8116ea,
32'h3d8c6554,
32'hbf562515,
32'hbfa8c902,
32'hbe6a3cdd,
32'h3dd1ca3e,
32'hbe286f3b,
32'hbe95fd44,
32'h3f064e01,
32'hbf116f31,
32'h3deaf947,
32'hbe91c823,
32'hbe6b5118,
32'hbe908034,
32'h3f11bda4,
32'hbef65280,
32'hbf185894,
32'h3eb158ad,
32'h3d8a9448,
32'h3ec2599b,
32'hbd8383d4,
32'hbe2a6d1e,
32'h3e73a922,
32'hbf88da00,
32'h3d48c0e2,
32'hbd509e8f,
32'hbdeed721,
32'hbf10bdb0,
32'hbda89c32,
32'h3da66653,
32'hbe9d8ea0,
32'hbe5b3692,
32'hbfa9c04a,
32'h3e5dc971,
32'h3ed4bd7d,
32'h3e0b847a,
32'hbee01daf,
32'h3e8fb500,
32'h3dad4531,
32'hbe5d7b52,
32'h3e2d64cf,
32'h3ca126b5,
32'hbebf10a8,
32'hbf5bb3ed,
32'hbe271e2a,
32'hbe19adbb,
32'hbd92f1c4,
32'h3d116e21,
32'h3dc42fe1,
32'h3ed3d696,
32'hbe11beff,
32'hbebdeac3,
32'h3d5c670f,
32'hbf37c155,
32'hbdccd58d,
32'hbcf2742a,
32'h3ee60fa1,
32'hbd8ad7ee,
32'h3d96a822,
32'h3d07bfbe,
32'h3d9e48db,
32'h3e60f77a,
32'hbf79b968,
32'hbf401a30,
32'hbf9933fe,
32'h3d06ab49,
32'hbed116fc,
32'h3cb44e50,
32'h3e7975d9,
32'hbf076599,
32'hbe6d58cf,
32'h3e8e7a80,
32'h3c5db5f2,
32'hbf3c1a8d,
32'hbe69d832,
32'hbf75b15f,
32'hbec17646,
32'hbccb8e57,
32'hbe449434,
32'h3eab8cb3,
32'h3e76d579,
32'h3dccfd56,
32'hbe022350,
32'hbf32ba39,
32'hbdf9c685,
32'hbd22da36,
32'h3d4890fb,
32'hbe8128ef,
32'h3d2eac4e,
32'h3e3c5960,
32'h3b5efde1,
32'hbd708d6e,
32'hbf211ca4,
32'hbf68c0d6,
32'hc016ed74,
32'h3e81409a,
32'hbeaf10e5,
32'hbe3167ad,
32'h3f0fbc6f,
32'hbbd67dbf,
32'h3e1a896c,
32'h3ed4f877,
32'h3d0f9c66,
32'hbf100a84,
32'hba854416,
32'hbfd464c4,
32'hbd97aa08,
32'h3c89f733,
32'hbe95ca9e,
32'hbdaa9e48,
32'h3dac95e8,
32'h3be68c1b,
32'hbe67227e,
32'h3f079ce5,
32'h3cc05cbb,
32'hbd9bb550,
32'hbe6471c2,
32'hbe698fbf,
32'hbde4242d,
32'hbd4f3211,
32'h3ee2584b,
32'hbeb88822,
32'hbf2c9f3f,
32'hbe6b3ccc,
32'hbe3a02f3,
32'h3decbb08,
32'hbe43731d,
32'hbe21571a,
32'h3dcce476,
32'hbf23a4be,
32'h3e36938b,
32'h3d923b7b,
32'hbe638094,
32'hbeb77aab,
32'hbe28457b,
32'hbf7b914a,
32'hbdbe7ba8,
32'hbd3121ec,
32'h3e4e594d,
32'hbd252dbb,
32'hbd06b93e,
32'hbe069650,
32'hbcd43aae,
32'hbe5c884d,
32'hbda7b7dc,
32'hbd4e3bf4,
32'hbeeec8cd,
32'hbddef605,
32'h3e169790,
32'hbd8823b3,
32'hbe9d82d9,
32'hbe7f7736,
32'hbf80a716,
32'hbe951faa,
32'h3f55cf6b,
32'h3e37e057,
32'hbdd701ba,
32'hbdb9b057,
32'hbd4141b8,
32'hbf2ff4fe,
32'h3df1415d,
32'h3d4eab36,
32'hbe498736,
32'h3de2d767,
32'hbdce7728,
32'h3e1089e6,
32'hbd374dfb,
32'h3dc3812f,
32'h3f006bb4,
32'h3de3c1d6,
32'hbd92fbc5,
32'hbd7925c3,
32'h3dcc0f03,
32'h3e8519a3,
32'hbd67c58c,
32'hbd322e9f,
32'hbe509307,
32'h3d907ddf,
32'h3e70661e,
32'hbe1abafe,
32'h3e1b9101,
32'hbe77a8db,
32'hbf68fbf9,
32'hbfa12053,
32'h3f141a13,
32'h3e1863e9,
32'hbd80ac13,
32'hbde6c22c,
32'hbd58e383,
32'hbe8de14c,
32'h3dfbc070,
32'h3aad994b,
32'hbbc2af1c,
32'hbe08b97a,
32'h3d968806,
32'hbdf3f40b,
32'h3e004096,
32'h3e8b83e3,
32'h3e588b73,
32'h3d7da0da,
32'hbd357bbd,
32'hbd9bbf6c,
32'h3dd3f2fa,
32'h3e4cbf07,
32'hbd6acec3,
32'hbb3afc1d,
32'h3ddfcfaf,
32'hbc9ed00c,
32'h3e4c3724,
32'hbd707871,
32'hbb953994,
32'hbe69cca4,
32'hbf23d380,
32'hbf8f9e23,
32'h3e8af7ea,
32'hbb6fae11,
32'hbdd1e024,
32'hbecc4097,
32'h3e810635,
32'h3e1cfd68,
32'h3e0a8e4a,
32'hbc766c8e,
32'h3e3b1932,
32'h3da3c17d,
32'hbe555124,
32'h3d59a9cd,
32'h3cf9f288,
32'h3ecbe932,
32'h3c53a529,
32'h3d8cc19b,
32'h3dbb5734,
32'hbe2f6a0d,
32'hbe39039a,
32'h3c993cf6,
32'hbdd773f5,
32'h3b9793d3,
32'hbcba677b,
32'hbd0b5323,
32'hbee0eb62,
32'hbe29198c,
32'hbe400197,
32'hbe017d4e,
32'hbef8ee81,
32'hbf1a790a,
32'h3e94b44a,
32'h3aaba0a8,
32'h3af71287,
32'hbca23a8b,
32'hbe7932ca,
32'hbd9b8c51,
32'hbdc30848,
32'h3e0ff45e,
32'hbe1746ab,
32'h3e6e2e59,
32'hbca40f3f,
32'hbd8d1a27,
32'h3dc2994e,
32'h3d4e45ee,
32'hbe858da2,
32'hbe00ed1d,
32'h3e213ba4,
32'hbc0b1571,
32'h3d74936d,
32'h3e32a84b,
32'hbc1a99c9,
32'hbd823ba5,
32'h3db6e4f2,
32'hbda1f3a7,
32'hbea42bad,
32'hbe7cfa54,
32'hbd108315,
32'h3dcaff2c,
32'hbe677915,
32'hbe1ab2a1,
32'hbdb2b08e,
32'hbdcd265b,
32'h3e51ef76,
32'hbea33e7c,
32'hbbb056b0,
32'hbeba0840,
32'hbe1199ff,
32'h3d1450f0,
32'hbe8bf052,
32'h3e9b6b0c,
32'hbe260622,
32'h3e0a7134,
32'h3b885811,
32'hbe29ffb2,
32'hbea4a547,
32'h3d698a82,
32'h3e1f65e6,
32'hbd8135d4,
32'hbdefac99,
32'h3e4d7d3d,
32'hbc8d9863,
32'hbc6afe84,
32'hbd8f6b44,
32'hbec86d67,
32'h3dc4b55f,
32'hbe01d4c7,
32'hbe02d0f1,
32'h3d2965a9,
32'hbea2b3f0,
32'hbd9c6509,
32'hbe407df4,
32'h3ed6e94e,
32'h3f03f6a8,
32'hbccebc25,
32'h3df43ba3,
32'hbe16aa3b,
32'h3d9e48b5,
32'h3d9d6f04,
32'hbef003d0,
32'h3e8bb2ab,
32'hbea4a45b,
32'hbd21064e,
32'h3dc95409,
32'hbbc659f5,
32'hbfafb366,
32'hbca5a175,
32'h3e3df9e1,
32'h3d5f7ce2,
32'hbe900b83,
32'hbdc29783,
32'hbdc78f15,
32'h3d33f736,
32'hbb41ec72,
32'hbeb7c8d2,
32'h3daf11c6,
32'hbdd6568f,
32'hbd9a2427,
32'h3d11bcfc,
32'hbeb2d148,
32'hbdd64e71,
32'hbe382334,
32'h3dc37a5c,
32'h3e937ee4,
32'h3c24eac5,
32'hb93868cb,
32'hbcce9031,
32'h3d8bfffa,
32'hbe2543d7,
32'hbf6974b9,
32'h3c3b4a5c,
32'hbef7118a,
32'hbea7b8cd,
32'hbd8ef883,
32'h3df32876,
32'hbf813447,
32'h3c2daad3,
32'hbcf004d9,
32'hbd4cfb2c,
32'hbe928bfb,
32'h3e5fb8f6,
32'hbd6f2d0f,
32'hbd3e4cdf,
32'hbd6d1e6a,
32'h3c95321a,
32'h3f03db5d,
32'hbd8f0441,
32'h3dcd83e6,
32'h3e8e11ab,
32'hbee8a7fc,
32'hbc593640,
32'hbe596486,
32'h3bf667aa,
32'h3ce86765,
32'hbe066c0c,
32'hbd412889,
32'hbe676bc5,
32'h3e1f76fc,
32'hbc98b8f0,
32'hbf3ba075,
32'h3e53b36f,
32'hbf26dda7,
32'h39832837,
32'hbca1d994,
32'hbe60c1f4,
32'hbfded06c,
32'h3e407750,
32'h3dfbbf43,
32'hbe26c02f,
32'hbebc36c8,
32'h3ea3d96e,
32'h3ae184fd,
32'h3dbb4664,
32'hbd0d6879,
32'h3cccdb0a,
32'h3e8d1928,
32'hbdcc9fed,
32'h3d1c13b0,
32'hbe6d6511,
32'hbe6712a2,
32'hbdf14d55,
32'hbd1b73d9,
32'hbc0b1590,
32'h3e2adad0,
32'hbc60577c,
32'hbe888e35,
32'hbd9464b4,
32'h3e3b7004,
32'h3e1cb9b9,
32'hbf6a51c5,
32'h3e2de42b,
32'h3dd33dda,
32'h3e43b461,
32'h3e60357c,
32'hbe22d41e,
32'hbfd2fd60,
32'h3e784cb2,
32'hbe9c5b24,
32'hbdd55a27,
32'hbf1a125b,
32'hbefbe0e1,
32'hbc88affb,
32'hbc95e7cb,
32'h3d6d2fd5,
32'hbe02ece4,
32'h3eb10a36,
32'h3e4849c4,
32'h3dadb073,
32'h3e4b32a2,
32'hbec0b627,
32'h3e7a106d,
32'hbe7f189e,
32'hbd4b8c49,
32'hbc999e0a,
32'hbb8a00f4,
32'hbe8fb9c6,
32'hbe80bdc0,
32'h3e132661,
32'hbdefe790,
32'hbf48c898,
32'h3e33b55a,
32'hbf3323c6,
32'h3d9f0197,
32'h3d540334,
32'hbea1759d,
32'hbde70482,
32'h3d9d787a,
32'hbd08086a,
32'hbdeea8d4,
32'h3e1bc17a,
32'h3e81a13a,
32'hbd70a914,
32'h3d19f069,
32'hbdd8c30c,
32'h3d60de87,
32'hbd7becf8,
32'h3e1e96c9,
32'h3d99643d,
32'hbc7496ca,
32'hbe93b63b,
32'h3e160656,
32'h3e103488,
32'h3dc55927,
32'hbc64897b,
32'hbdcd78bb,
32'hbdcb2f1c,
32'hbf3bad49,
32'h3e45afb5,
32'hbe1869f1,
32'hbe38e4b7,
32'hbbc4de2f,
32'h3d904084,
32'h3d21c570,
32'h3d619a5a,
32'hbeddfda8,
32'hbe558455,
32'hbdf18921,
32'hbda31db4,
32'hbddc26a9,
32'hbee1a7ad,
32'h3d06b10e,
32'hbdfc8a48,
32'hbd3a0544,
32'hbf020ba5,
32'h3ebb5c80,
32'h3d8a22c1,
32'h3cf6b2ec,
32'h3ef7de92,
32'hbdd4f379,
32'hbf1b2bfc,
32'hbe037f9b,
32'hbd0350ac,
32'hbdb9b407,
32'h3e1347d8,
32'hbd8c0766,
32'hbe3c3d02,
32'hbf7e7cb5,
32'h3e3c584e,
32'h3dd431ae,
32'h3e48a77e,
32'h3e967219,
32'hbf5d997c,
32'hbe772423,
32'hbb91d258,
32'hbea7bddc,
32'h3ed9d059,
32'hbdd82d13,
32'hbe32ec69,
32'hbe7f6cb5,
32'hbe62f62e,
32'h3e7c5dcc,
32'h3dfdda93,
32'hbd97c4ce,
32'hbf182b9c,
32'h3ec70cad,
32'h3e1f43c3,
32'hbd430847,
32'h3e5030f6,
32'h3f0ef33d,
32'hbf0f50e7,
32'h3edce3fa,
32'hbe3d23a1,
32'h3df5be19,
32'h3e9ba8fb,
32'hbc30eec5,
32'h3de2bfdb,
32'hbf771254,
32'h3df83c82,
32'h3df48639,
32'hbd01e62f,
32'hbf1ab396,
32'hbd4ea5f3,
32'hbcd74f30,
32'hbde9e154,
32'hbee68a17,
32'h3e96fbe2,
32'h3e2649d5,
32'hbed89e9c,
32'h3d859dac,
32'hbe97521b,
32'h3e6a78c2,
32'h3bc42527,
32'h3d39948b,
32'hbeda1b71,
32'h3f2be779,
32'h3d814b5d,
32'hbdb8f4aa,
32'hbd35ba88,
32'hbe4da603,
32'hbef9f8d7,
32'h3ea3ac53,
32'hbf061fd5,
32'h3e180118,
32'hbe007845,
32'h3e3b6ec0,
32'h3cea1644,
32'hbd350533,
32'hbda64132,
32'hbe2bcacc,
32'h3e60b5c0,
32'hbf82273d,
32'h3edef930,
32'h3e16de16,
32'h3ec5ff68,
32'hbe6eb26c,
32'hbde595da,
32'hbf44afbd,
32'hbe9dc302,
32'hbe99b315,
32'hbf342ce2,
32'hbe18ca47,
32'hbd8d5a11,
32'hbd0a997b,
32'h3e160b2a,
32'h3f181a97,
32'hbe000420,
32'hbe292a88,
32'h3f7e54ad,
32'h3e9c0d15,
32'hbf11589f,
32'hbba66dc2,
32'h3cf7c04c,
32'h3d1c0d66,
32'hbe13d9d2,
32'h3e2caa56,
32'hbdce6961,
32'hbe88e431,
32'h3e68f861,
32'hbd0c85dc,
32'h3eb34127,
32'hbf62ddad,
32'h3ed8544e,
32'hbeb9e4f2,
32'h3f4d9dff,
32'hbd10f904,
32'hbd8d7352,
32'hbf8c0654,
32'hbe30fb5f,
32'hbebb3b48,
32'hbf1bc46b,
32'h3d1fc8e6,
32'h3ae5a30b,
32'h3defb9d5,
32'hbefaca70,
32'h3ec2134f,
32'hbe63853c,
32'hbecfb486,
32'h3dede45f,
32'hbe1362ae,
32'hbf83fb41,
32'h3edfd493,
32'h3c1087ee,
32'h3ebc3fc0,
32'h3eeb8ea1,
32'hbec20f7f,
32'hbe80a089,
32'hbf352f60,
32'h3f21507b,
32'h3f0b41f2,
32'hbdbdccc5,
32'hbe90fbfd,
32'h3ee678cf,
32'h3f28d359,
32'h3ebd4b84,
32'hbdaf9317,
32'h3ec003ba,
32'hbe239ea0,
32'hbf10a6e1,
32'hbef9b107,
32'hbebf808f,
32'h3e2f8414,
32'h3c4c366d,
32'h3d763265,
32'hbf429785,
32'h3f1afd50,
32'h3f1c479f,
32'hbe8077db,
32'h3f1ecfcd,
32'h3e99f171,
32'h3f059be1,
32'h3f49844b,
32'hbefdc9ac,
32'hbb8fe9e5,
32'hbfaad0a8,
32'hbee961a0,
32'h3ef691a6,
32'hbd8a774f,
32'h3e97754c,
32'hbe3f6b10,
32'h3e9729fe,
32'hbf65c807,
32'h3f3565a0,
32'hbe203007,
32'h402fb347,
32'hbe49d9d3,
32'hbdbabca6,
32'hbe2704f4,
32'h3f156f15,
32'hbe8d880d,
32'h3e839f9c,
32'h3f7e99a3,
32'hbd003ded,
32'h3d76b496,
32'h3d273511,
32'h3f147030,
32'h3f695fe4,
32'hbf8affa6,
32'h3fdb33a5,
32'hbe8db88e,
32'h3f4c4868,
32'h3e4b0db8,
32'hbe8be12c,
32'h3d622a17,
32'hbec342e2,
32'h3e3bee48,
32'h3f69e725,
32'h3d3884bb,
32'h3ed9c08f,
32'hbf381f8f,
32'h3ed588e0,
32'hbf2a7d0b,
32'h3f662493,
32'h3d831bed,
32'h3f9387e3,
32'h3fcd7a68,
32'h3b690bc2,
32'h3eee0d1d,
32'hbc873233,
32'hbee8af26,
32'h3eab2248,
32'h3f346be0,
32'h3d2a73b7,
32'hb9de660d,
32'h3f436cab,
32'hbeeff227,
32'h3e2a019a,
32'hbf3b0e8f,
32'h3f929b02,
32'h3d20f4fc,
32'hbf920753,
32'hbed5e3b5,
32'h3b8c262f,
32'h3f386982,
32'hbdbe2270,
32'h3efccaf2,
32'h3ec059f2,
32'h3d889df2,
32'h3e13a3b0,
32'hbeba62d3,
32'hbe055134,
32'h3ee62f97,
32'h3de60b6c,
32'hbdbc712d,
32'hbd49b8ed,
32'hbd660ba8,
32'h3db30ba6,
32'hbd4455be,
32'hbd96f3bb,
32'hbd5b2d93,
32'h3d0dab56,
32'h3d2f6041,
32'h3ce68d3e,
32'hbd4f1340,
32'h3cdbeefc,
32'h3c1cff66,
32'hbd3e4df1,
32'h3d095c04,
32'h3bada282,
32'hbbb92ddf,
32'h3cb21432,
32'h3d0c4721,
32'hbda36779,
32'h3c6c6dcc,
32'hbc9411f3,
32'h3c085c42,
32'hbce5e981,
32'h3d641a66,
32'hbd9c97ba,
32'h3d910ad4,
32'h3d1b302b,
32'h3ad93a5a,
32'hbcf5ccdf,
32'h3d90c007,
32'h3d327d84,
32'hbd9edd9c,
32'h3d9e563a,
32'hbd6334b9,
32'h3d94f37b,
32'h3d0a2284,
32'h3d8171be,
32'h3dd3a9c8,
32'h3dbeaa96,
32'h3c8561e6,
32'h3dccec6d,
32'hbbba2bfd,
32'h3be39fb7,
32'h3dd14d4b,
32'hbd918b6e,
32'h3b5f9d68,
32'h3c46cefd,
32'hbc93cfeb,
32'h3db9e8a2,
32'h3db23456,
32'hbdab82c9,
32'hbca3eb9f,
32'hbcc6c946,
32'hbc15a75b,
32'h3c1fdd7b,
32'h3c8dbb6f,
32'hbd88854f,
32'h3d32f6a3,
32'hbd8123c2,
32'h3dc991c2,
32'h3da13b20,
32'hbd345381,
32'h3b983269,
32'hbdedb025,
32'h3e83b62a,
32'h3c56c5ac,
32'h3cc2e1b4,
32'h3cce6e07,
32'hbd9e3938,
32'hbd9d359f,
32'hbc01ad8c,
32'hbddf1425,
32'h3dc60a8d,
32'h3e5a55c3,
32'h3d52b853,
32'h3d8750bc,
32'h3ccf78a9,
32'hbc00c536,
32'h3d4fb772,
32'h3edc90fe,
32'h3cb1969b,
32'hbd9fde4b,
32'h3e82e086,
32'h3d5dccb7,
32'h3e122f0b,
32'hbd8dc055,
32'h3c615fa6,
32'h3d710067,
32'h3e0097a7,
32'h3e402390,
32'h3fc0ecb9,
32'h3d5c916e,
32'hbdfa8e66,
32'hbd978816,
32'hbd87be2c,
32'hbe6cb3c3,
32'h3eb4a04c,
32'h3affb0eb,
32'h3b827b09,
32'h3cd5e6dd,
32'hbec12346,
32'h3f2c33da,
32'h3ed9c0cf,
32'hbe1056cd,
32'hbe3b7a47,
32'h3e0da9e7,
32'hbe4b9704,
32'hbe8c5e16,
32'hbdbc5705,
32'h3ee70e83,
32'hbc7cb11f,
32'hbd6b65b4,
32'hbb61f6cc,
32'hbd332bdb,
32'hbe819bfe,
32'h3f0a5c7e,
32'hbeb98a8e,
32'hbe001e2e,
32'hbdf48563,
32'hbf5ecec7,
32'h3ea719a2,
32'h3de31120,
32'h3eda50d6,
32'h3e0a19b7,
32'hbe00fd2f,
32'hbdad5225,
32'h3e6ea7fd,
32'hbda87581,
32'hbdbc8ca2,
32'hbdb44ea8,
32'h3e6bbce5,
32'h3f8a038b,
32'h3d0e3ba3,
32'hbeebe42d,
32'h3fa55409,
32'hbea941dd,
32'hbec22d47,
32'hbfc51c42,
32'hbee98f7c,
32'h3df7bc2b,
32'hbbcb04ff,
32'h3bad6afa,
32'h3e04ab67,
32'hbf0b88de,
32'h3de78730,
32'hbee55d95,
32'h3cee765c,
32'hbe6a1a4c,
32'h3f546521,
32'hbf4e99aa,
32'h3dc60cad,
32'hbec13af7,
32'h3f1c8ef6,
32'hbee13a16,
32'h3e4d4319,
32'hbdebbd31,
32'h3e97d011,
32'hbe1e9850,
32'hbbcf9a21,
32'hbd834509,
32'hbe9ed27b,
32'hbe6f147b,
32'h3bda0099,
32'h3d5c2da9,
32'h3db8f8e5,
32'h3f4b004b,
32'hbfa8e6b8,
32'hbfd3fd83,
32'h3e3b9136,
32'hbda3b1f5,
32'hbe06c377,
32'h3ecc7292,
32'hbe31c266,
32'hbeb10065,
32'h3cc2afcd,
32'h3e87768f,
32'hbeb5a5d7,
32'hbfd00a45,
32'h3eee1070,
32'hbe19e444,
32'hbf2257f9,
32'h3f38e541,
32'hbe1fe340,
32'h3ed3bbfd,
32'h3d132264,
32'hbeb56021,
32'h3d5d3a7e,
32'hbee8dec0,
32'hbd025a7d,
32'hbd95e588,
32'h3d6bc644,
32'hbe837c09,
32'h3e900c52,
32'h3e604ad2,
32'hbe05aa91,
32'h3ed03d00,
32'hbfa4c513,
32'hbe58997d,
32'hbf540e08,
32'hbca1531c,
32'hbf2e4910,
32'hbea062ed,
32'h3e64dff9,
32'h3d69f23e,
32'hbd018f91,
32'h3e5cccb5,
32'h3e4e402f,
32'hbfbc33c9,
32'h3daecbe2,
32'hbf7227e2,
32'hbe96f37a,
32'h3db18ed3,
32'hbd772d9e,
32'hbe763b26,
32'h3ec5f5bc,
32'hbefe9f7b,
32'h3deffd61,
32'h3d04db8b,
32'hbb8f20bf,
32'h3c841c65,
32'h3f1622f9,
32'hbe39bc71,
32'h3e46cff1,
32'h3eb123a0,
32'h3e4a9c8e,
32'h3dacc047,
32'hbf81efc2,
32'hbf5ec5fc,
32'hbe691f86,
32'h3ca787ec,
32'hbfe0dc89,
32'h3de71437,
32'hbebb5f12,
32'hbced3900,
32'hbe046818,
32'h3c9b84af,
32'h3ea1fb09,
32'hbf8d99d0,
32'hbe128785,
32'hbe0e285d,
32'h3e07f434,
32'h3e3d75f3,
32'h3e5feefd,
32'h3d1560ca,
32'h3eabf68e,
32'hbe0e1448,
32'hbdc227a1,
32'h3e75c0aa,
32'hbd1f843d,
32'hbc913c18,
32'h3e86a448,
32'hbe79e1fc,
32'h3d169be5,
32'h3e5e227a,
32'h3e1d1ed6,
32'hbe0f0aab,
32'hbfa1a3ea,
32'hbfa905ea,
32'hbefe7bf2,
32'hbe3063f2,
32'hbe3509c6,
32'h3e0988e6,
32'hbafd7c96,
32'h3de932b6,
32'hbe5c9563,
32'hbef03fc0,
32'h3d92cb90,
32'hbf9955f3,
32'h3e15a86d,
32'h3ee665f0,
32'h3e257710,
32'h3e3f882f,
32'h3e17d83c,
32'hbd8027ba,
32'hbe4db0a1,
32'hbe761922,
32'hbd30b9ac,
32'h3e2d95f8,
32'h3aeb000c,
32'hbd23c08e,
32'h3cfa5d04,
32'hbe536027,
32'h3eabb1a7,
32'h3ce45f6b,
32'h3d5202e9,
32'hbe6847e9,
32'hbe028649,
32'hbfd885cc,
32'hbe2f1279,
32'h3e113608,
32'hbe9d6571,
32'hbe5c45ad,
32'h3d658db5,
32'h3e3156eb,
32'hbd8926a8,
32'hbd96c55c,
32'h3e54235d,
32'hbe9941fc,
32'hbd46cc8f,
32'h3e90565a,
32'hbd2b1d66,
32'h3ceeeb23,
32'h3e1ee238,
32'hbdd87653,
32'h3d674e73,
32'hbe02523e,
32'h3ce124f6,
32'hbdb672c6,
32'hbd67ea15,
32'h3da1ac33,
32'h3e009aad,
32'h3d48438d,
32'h3e6af2c3,
32'h3d81bc8c,
32'hbdb55d3a,
32'hbd9d0482,
32'h3ce8445b,
32'hbfcd6688,
32'hbe467771,
32'h3eb82721,
32'h3d9c796c,
32'hbe8ff953,
32'hbe284dda,
32'h3e960301,
32'h3e384ae5,
32'h3daa0c3e,
32'hbdc2ad11,
32'h3d453a6b,
32'hbe3670b4,
32'hbe821709,
32'h3d85de9c,
32'h3e4fc1b4,
32'h3d6be625,
32'hbebd58f4,
32'h3df427bf,
32'h3cacdf86,
32'hbefaf0fa,
32'h3e4b58b4,
32'h3cf1a4c8,
32'hbd8087b6,
32'h3ebb29c8,
32'h3eb02bac,
32'hbe353f94,
32'hbe5f3141,
32'hbec2a681,
32'hbe3dce4a,
32'h3d99defb,
32'hbf0195b6,
32'hbe5084e3,
32'hbbddd1d8,
32'h3debcf42,
32'hbe67bfc0,
32'h3b6b82d8,
32'h3e418732,
32'h3e01ad6b,
32'h3d2e793f,
32'hbd56df9c,
32'hbe579311,
32'hbeb3a6e9,
32'hbe1ec2fc,
32'h3eae37a5,
32'h3e22c126,
32'hbd7d6316,
32'hbea44982,
32'h3d3644b9,
32'h3cd322a9,
32'hbe8b6f13,
32'hbeb9473b,
32'hbd036998,
32'hbd484056,
32'h3eb8e4c3,
32'h3e645f12,
32'hbe2e9ac6,
32'hbe64ea52,
32'hbbbd986a,
32'h3cf9588a,
32'hbec183cf,
32'hbcf126d0,
32'hbe923c84,
32'h3dce316d,
32'hbe887a8c,
32'h3b99ad8f,
32'hbd33bf7b,
32'h3d212acd,
32'h3e9504c2,
32'h3dc0a3f4,
32'hbcc23be8,
32'hbd8a5c5b,
32'hbef397f2,
32'hbd05fbd4,
32'hbd391aa6,
32'hbcea1d03,
32'hbca65b03,
32'hbdc6680b,
32'hbe3c38e4,
32'hbe38aec2,
32'h3e241b90,
32'hbd992cb2,
32'hbd8ddbeb,
32'hbce1e3ee,
32'h3b219830,
32'h3d0ef0b1,
32'hbe25c792,
32'hbd0998c5,
32'hbe8e2503,
32'h3c81f609,
32'hbecbcb87,
32'h3bb44ab2,
32'hbe9d97e7,
32'hbcacdaf7,
32'h3e1a7376,
32'hbe074a43,
32'hbe824bcb,
32'hbe5e7278,
32'h3e4bce40,
32'hbc92982a,
32'h3e36193c,
32'h3e460e99,
32'h3cd94723,
32'hbd9640e4,
32'h3e325f80,
32'h3cba0fad,
32'hbee05936,
32'hbd8b45e0,
32'hbddc3b2b,
32'hbe801a59,
32'hbeb01a83,
32'hbdded840,
32'h3c5d8508,
32'hbd821fab,
32'hbe91474c,
32'hbe76a563,
32'hbe204ce4,
32'hbe0c6f51,
32'hbd960feb,
32'hbd6cb9f6,
32'hbea49698,
32'hbe5a7ffe,
32'hbee6658c,
32'hbd0b1145,
32'h3e444761,
32'h3d277902,
32'hbccb544e,
32'h3d8179e1,
32'h3e3a9f6a,
32'hbca76002,
32'hbece0292,
32'hbd402f88,
32'h3e65e2b4,
32'h3e20ee26,
32'h3dee93aa,
32'h3d861f60,
32'hbfdbc430,
32'hbd10d461,
32'hbdb3b5f0,
32'hbeb2e122,
32'hbd8fb765,
32'hbe29438e,
32'h3ca7d3d5,
32'h3c97d383,
32'hbeb2dafe,
32'hbef325f5,
32'hbec7eaad,
32'hbe3fd12e,
32'h3eedd08c,
32'hbe0ebc72,
32'hbe9a9f8f,
32'hbe344ae6,
32'hbe84b6c6,
32'hbd3555a7,
32'hbd870f11,
32'hba9f0cd8,
32'hbe4ed8db,
32'hbeb10892,
32'h3df0be04,
32'h3b86a584,
32'hbf8fc315,
32'h3bd43218,
32'hbf0d1a7b,
32'h3da2c306,
32'hbe10927e,
32'hbd7a4a48,
32'hbe14accd,
32'hbe07f166,
32'h3d531c08,
32'hbcb6774b,
32'hbe9ca4aa,
32'h3c8859bc,
32'h3d599bc3,
32'hbc5aee6e,
32'hbf09136d,
32'hbf0262a8,
32'h3d70de27,
32'hbe3442d5,
32'h3e8810fa,
32'hbc9c35cb,
32'hbe72c49e,
32'hbe2e87d6,
32'hbe00c1dd,
32'hbe2ede4e,
32'h3e291dc1,
32'hbe1087ff,
32'h3dc9690d,
32'h3e580da1,
32'h3d790f24,
32'hbe33cbc3,
32'hbf283d22,
32'h3e8078dc,
32'h3e662e28,
32'h3cf296ba,
32'hbead6335,
32'hbc2309a4,
32'hbe9c2c31,
32'h3d136654,
32'h3db7c4e5,
32'hbdb8ac23,
32'hbf5bd6f9,
32'h3dfac799,
32'hbd5f8e9d,
32'hbdf99d64,
32'hbd5c52a4,
32'hbeec7787,
32'h3e0725a0,
32'hbe4c2e05,
32'h3ed411f0,
32'hbe4f5d56,
32'hbe80216f,
32'hbed7b649,
32'h3ed3f576,
32'h3c93db95,
32'h3df46a0c,
32'h3bf530fb,
32'h3e21a971,
32'hbca647ab,
32'hbd278791,
32'hbe31bce0,
32'hbf240ab1,
32'h3e6510d7,
32'hbefdf283,
32'h3e9b1929,
32'hbc25bcc0,
32'h3e4d1f8c,
32'hbea6eacf,
32'h3db6a7d0,
32'hbe1dc135,
32'h3e94bffb,
32'hbf5d1f20,
32'hbea1427b,
32'hbd3866fb,
32'hbcf419ef,
32'hbd954338,
32'hbdb5e774,
32'h3ee291f5,
32'hbe50dd5d,
32'h3ecf7668,
32'hbe1fcf2c,
32'hbe656e5d,
32'hbe3799a8,
32'hbdea4df6,
32'h3da664f1,
32'h3d2c8a57,
32'h3ddb5406,
32'h3dbe18fa,
32'h3e11f235,
32'h3d8fa91f,
32'hbd8248df,
32'hbf50e4ae,
32'hbe26e429,
32'hbf7fc064,
32'h3e8f0042,
32'hbd2a01a2,
32'h3e89f70d,
32'h3f2c425c,
32'h3e822fdb,
32'h3dd6bb71,
32'hbe312943,
32'hbeb6aee9,
32'h3efca877,
32'hbd6cd52e,
32'hbdaa82f6,
32'hbd1ce279,
32'hbe1fce30,
32'h3ec68172,
32'hbd52142e,
32'h3f472858,
32'hbed7816f,
32'hbe806551,
32'hbe013659,
32'hbe24f9d6,
32'hbdebccf1,
32'hbeef1d67,
32'hbe096f1b,
32'hbed52ca1,
32'hbeb9ae20,
32'h3e56f2cd,
32'h3e06efe4,
32'hbeb05a33,
32'hbd9eb183,
32'hbe170434,
32'h3e9aab3d,
32'h3eef4d4b,
32'hbd4a966f,
32'h3e69c71c,
32'h3e3c4c58,
32'h3e63ea6d,
32'hbed5cdf3,
32'hbfab6bbf,
32'hbe05bcc7,
32'h3cd7a759,
32'h3d01a951,
32'hbf0d29fc,
32'h3d95a373,
32'h3e1d14fa,
32'hbd9cb103,
32'h3efda91d,
32'hbd8deced,
32'hbdca0e82,
32'hbe18c395,
32'h3f07aa3b,
32'hbefc48bb,
32'hbed8ee76,
32'hbe10d321,
32'h3e825a4a,
32'hbf3cab3e,
32'h3ddfbca2,
32'hbe27292f,
32'hbe4cd722,
32'h3df3a652,
32'hbee60996,
32'h3e248e47,
32'hbc4b55f2,
32'h3ea78f7d,
32'h3f099bae,
32'h3e89391d,
32'h3d34e480,
32'hbe32e48b,
32'hbf7b4d3e,
32'hbd605747,
32'h3ca0f740,
32'hbc4b3006,
32'hbe43da72,
32'h3df2c7f2,
32'hbe040ed1,
32'h3dc32d97,
32'hbeb97d33,
32'hbe851ef2,
32'hbe553372,
32'hbe6b5333,
32'h3eadc5db,
32'hbd5b56ac,
32'h3e443699,
32'hbe216dc5,
32'h3da0bd06,
32'hbedfbf4a,
32'h3e59a3ce,
32'h3e2c8ef1,
32'hbf05f2b0,
32'hbf0f1d53,
32'hbdb9a6fa,
32'hbd77c0fe,
32'h3ec82ecb,
32'hbe87b23e,
32'h3eb76777,
32'hbcbead97,
32'hbea9786f,
32'hbf817fba,
32'hbf617ee9,
32'h3e339556,
32'h3d66d93d,
32'h3ca69583,
32'hbe2ced5f,
32'h3e408559,
32'h3ec1f135,
32'h3c0fa3f0,
32'h3d4eea8e,
32'hbdeb4bff,
32'hbee1899f,
32'h3cfeb765,
32'h3db5b05d,
32'hbd4da513,
32'hbf2ea57d,
32'h3e85368d,
32'hbe82bfda,
32'hbe7f36dc,
32'hbd9e47d8,
32'h3e20620c,
32'hbf25208d,
32'hbda3abf7,
32'h3ebe653a,
32'hbe94440f,
32'h3e794d5b,
32'h3d51712c,
32'h3d80ae1c,
32'hbf124d28,
32'h3cb6a955,
32'hbf84ed1a,
32'hbf57b0c6,
32'h3d37e57e,
32'h3ba5fc02,
32'h3d10c01d,
32'hbd923be4,
32'h3ed2f8d9,
32'h3e04d952,
32'hbe7cd7d3,
32'h3e9034ac,
32'h3dce01e0,
32'hbe500fab,
32'h3e462f8f,
32'hbe774d99,
32'h3e051392,
32'hbe6b6a83,
32'hbef6cce0,
32'h3b4405dd,
32'hbef8d83e,
32'h3ef5275d,
32'h3e44e12f,
32'hbdc6effc,
32'hbdaabca2,
32'h3edf40ed,
32'h3d138c9c,
32'h3e2e24d4,
32'hbf156d93,
32'h3eb7dfc3,
32'hbe9802d3,
32'h3f57672c,
32'h3edb6b4a,
32'h3db40fc3,
32'h3f01918e,
32'h3d1a8ae2,
32'h3c19cded,
32'hbf89b554,
32'hbdcb5b8f,
32'hbd54a02e,
32'hbd000b2c,
32'hbedff578,
32'hbf3c47aa,
32'hbd8a312d,
32'h3d05121a,
32'hbf70d8be,
32'h3e6508ec,
32'hbe3af2aa,
32'hbe7b50c6,
32'h3e8a739f,
32'hbf538b08,
32'h3f81b647,
32'h3df5e479,
32'hbdaf72e7,
32'hbf97cf59,
32'h3ee93621,
32'hbcd1bc67,
32'h3e564701,
32'hbf5fb237,
32'hbdef873e,
32'hbf086945,
32'hbe8652fb,
32'hbf2ff727,
32'hbd6e3ac5,
32'h3f44e2f5,
32'h3d669359,
32'hbc80d60d,
32'hbf483338,
32'h3ee6226b,
32'h3ef40f4d,
32'h3df32f3a,
32'h3f67b6e6,
32'hbe9fb400,
32'h3daf6062,
32'hbe10900e,
32'hbf4502c1,
32'h3e30c5c1,
32'hbf4fc072,
32'h3f5419e4,
32'hbe2b9cf1,
32'hbc3e8e14,
32'h3efc4dd1,
32'hbec1e526,
32'h3ec5fb86,
32'hbeb20fbb,
32'h3cf19eef,
32'hbd4595d3,
32'h3f48bf13,
32'h3e1083b8,
32'hbe390805,
32'hbe00ba9b,
32'hbde27c8b,
32'hbe73d5e4,
32'h3f08f270,
32'h3fa333be,
32'hbd9b3ebe,
32'h3d90c629,
32'h3f3c922e,
32'hbf06cac9,
32'h3ecb7e59,
32'hbe776e58,
32'h3fcb7ce5,
32'h3e0583ec,
32'h39aa3148,
32'hbe4f8d69,
32'hbf11280e,
32'h3c9eb106,
32'hbf27f825,
32'h3f691ad4,
32'hbd86d1b0,
32'h3ec52e79,
32'h3e57d45a,
32'hbf3c13f6,
32'h3f2bedfa,
32'hbeb6d1bd,
32'h3f542ff6,
32'h3ddea3cd,
32'h3dede7e4,
32'h3fec2dac,
32'h3d492a0a,
32'h3e5c67e7,
32'hbeff0d25,
32'h3d8abcfb,
32'hbd810a01,
32'h3f79a387,
32'h3d1496b0,
32'hbda92022,
32'h3fb3c61f,
32'hbfa2219e,
32'h3c106725,
32'hbf7c2efb,
32'h3eacd3b7,
32'h3f4a9f6c,
32'hbf9661ae,
32'h3ed231bc,
32'h3f26bc22,
32'h3ed33157,
32'hbe256e23,
32'h3f5d2b01,
32'h3e45cf30,
32'h3d8d92ed,
32'hbf2cfe8a,
32'h3d932d24,
32'hbf2409d6,
32'h3f67f8e8,
32'h3bb9fcd4,
32'hbbd8acc4,
32'h3c285d52,
32'hbd27856a,
32'hbc9bbda2,
32'hbbfe344e,
32'h3da1f267,
32'h3c89e1e6,
32'hbdba136c,
32'hbcdb7294,
32'h3dae56e2,
32'hbd31be11,
32'h3dc312da,
32'h3cf666d9,
32'hbd6d5c6a,
32'hbd848165,
32'h3d156f3a,
32'h3cdf2feb,
32'h3d4aac9e,
32'h3ddd9885,
32'h3cefb4a4,
32'hbdf7f5d0,
32'hbb86fd56,
32'hbd9a64ca,
32'h3d6e0a16,
32'h3ccf1e13,
32'h3cdd0ba3,
32'h3d8a546d,
32'hbd08e9b1,
32'hbcc5e574,
32'h3ceb36a5,
32'h3d8e6712,
32'hbd964715,
32'h3d4ef309,
32'hbd461c13,
32'h3d995530,
32'h3cab0fba,
32'hbd4593ea,
32'h3dbb548e,
32'hbd68177c,
32'h3d9a0801,
32'h3bd11297,
32'hbc984228,
32'hbd040978,
32'h3c4c0cee,
32'hbc016708,
32'hbcd4d164,
32'h3d043565,
32'h3caa09d5,
32'hbd3d7822,
32'h3cbb0a77,
32'h3cf7e208,
32'h3d849cc5,
32'h3c8b3f78,
32'hbd8cf870,
32'hbdb48d14,
32'h3b840c84,
32'h3c2497ab,
32'h3d7e06fd,
32'hbdea4faa,
32'h3c8af14c,
32'h3ca08b72,
32'hbc8b70ca,
32'hbd4255c7,
32'hbd587600,
32'hbd2f2a71,
32'hbdc5a209,
32'hbd3eeabf,
32'h3cee9444,
32'hbddecc6b,
32'h3d44a876,
32'h3cb7f00c,
32'hbab8ab59,
32'hbd90ad03,
32'h3bdbfff1,
32'h3cb5d622,
32'h3cb5ec5d,
32'h3d456dc8,
32'h3d91d1d7,
32'hbd81b704,
32'hbd8b3d1f,
32'hbd16b9f6,
32'hbb4bf5b1,
32'hbd7c1f11,
32'h3c42d0fc,
32'hbcf22d00,
32'h3d62578f,
32'hbd34d5c1,
32'h3ca5818f,
32'h3d48ccff,
32'hbe145229,
32'h3ec968e1,
32'h3f202bcf,
32'hbe0835e3,
32'hbec14c7f,
32'hbe864568,
32'h3eb9e0d9,
32'hbee03bfd,
32'h3e3c5739,
32'hbd32be96,
32'h3d81b6c0,
32'hbd051992,
32'hbecb0567,
32'h3f1c8a63,
32'h3eb2f528,
32'hbe4c5e4b,
32'h3bc96552,
32'h3d40f380,
32'h3c845912,
32'hbd30df02,
32'hbe7195ca,
32'h3ca58d68,
32'hbdc8d1fe,
32'hbf0262ca,
32'h3ee3de12,
32'hbdd02196,
32'h3f3415bb,
32'h3f3d1fff,
32'hbea81c51,
32'hbe665cae,
32'hbf7bc210,
32'h3eb208dd,
32'hbeab3552,
32'hbf4868b6,
32'hbe879a95,
32'hbf55a2d6,
32'h3ee7c44a,
32'hbe8e437e,
32'hbe8ef276,
32'hbc7b3d09,
32'h3d71a17e,
32'hbddb5b0d,
32'hbf5113dd,
32'hbf207469,
32'hbe7fe2d5,
32'hbe827489,
32'h3f9ecd06,
32'hbf373db1,
32'h3c954e6e,
32'hbed7b271,
32'hbf0e857e,
32'h3e8e6535,
32'hbdc1dc9e,
32'h3e2942d7,
32'hbea23436,
32'hbf54fded,
32'h3ed0c03a,
32'hbd7b86a0,
32'h3eb78da2,
32'h3e7f40e6,
32'h3e2fccf7,
32'h3f0dd08f,
32'hbf04748f,
32'hbf96a79f,
32'hbd65bba8,
32'hbf19f690,
32'h3e8dfed2,
32'h3e50888e,
32'hbd825f74,
32'hbf36befb,
32'hbb7ab1d9,
32'hbc86abb9,
32'hbf506d57,
32'hbe33e8a5,
32'hbe35b0fc,
32'hbd160805,
32'h3e2143e9,
32'hbf453aad,
32'hbfa738d0,
32'hbf886484,
32'hbfa85c57,
32'h3f252679,
32'hbcbf8a94,
32'h3ef88eb4,
32'h3f14f4ae,
32'hbd8fac9f,
32'h3f47a68b,
32'h3f444cb4,
32'h3cc5b2ab,
32'hbe92aa96,
32'h3f0eb12f,
32'h3ed4359e,
32'h3ded8290,
32'h3ed1345f,
32'hbe299b49,
32'h3f1e8dd9,
32'h3e803e9e,
32'h3d2d49b7,
32'h3d8a2697,
32'hbf717e12,
32'hbd2886cb,
32'hbcf70d02,
32'hbdbb3221,
32'h3eb800ca,
32'h3eaa776e,
32'hbdc3c52b,
32'h3d80678a,
32'hbf13cb8f,
32'hbf2563b8,
32'hbf038cc0,
32'hbf490745,
32'hbdde477c,
32'hbeadde05,
32'hbee7728a,
32'h3f3128b8,
32'h3f805da3,
32'h3f59639e,
32'h3effdaae,
32'hbb165a54,
32'hbee83031,
32'h3e61a45f,
32'h3ef8b256,
32'h3ef5ece2,
32'h3e6d6504,
32'h3ec2fac3,
32'h3e4940af,
32'h3e61a6ab,
32'hbec661d2,
32'hbdcd3e56,
32'hbdf3f895,
32'hbcd8f2ae,
32'h3c73a75d,
32'hbe1a3d5a,
32'hbe5d8bd5,
32'h3e975b07,
32'hbd92c3f3,
32'hbe32cfd6,
32'hbe972c52,
32'hbebcc4ce,
32'hbf07208d,
32'hbcfb4b20,
32'h3c9dfa2f,
32'hbf394dc8,
32'hbd1e7ce9,
32'h3e8ff08b,
32'h3f702dd9,
32'h3f039273,
32'h3be1390b,
32'hbc55dd92,
32'hbf5fc4af,
32'hbe8d497b,
32'h3ededbf7,
32'h3efc4277,
32'h3da767b9,
32'h3f2b2849,
32'h3dd8a594,
32'h3dd05f72,
32'h3cc49722,
32'hbeac1f6b,
32'hbf4d924b,
32'hbbd2658e,
32'hbdac8a82,
32'h3eb620bd,
32'h3d3ad6ed,
32'h3e813bb9,
32'hbdb4ad93,
32'hbe391dd8,
32'hbc42e663,
32'hbeb23d9b,
32'hbf5d3647,
32'hbec3dcb0,
32'h3e4c3ba5,
32'hbfaf4ff4,
32'hbc4a1a21,
32'h3d4f0e28,
32'h3f365a1e,
32'h3ec972f9,
32'hbbbafa2d,
32'hbeabc933,
32'hbe18b545,
32'h3e8f0938,
32'h3ded2781,
32'h3e1ef71e,
32'h3e5f9a66,
32'hbd6c28de,
32'hbd5ed606,
32'hba87094a,
32'h3e359ef0,
32'hbb546168,
32'hbd6a8602,
32'hbcf4210d,
32'hbd4962b8,
32'hbd0b05f3,
32'hbe871a6f,
32'h3e1c5576,
32'h3d4415d0,
32'h3e2fb35a,
32'hbd2b1e1d,
32'h3d84df9c,
32'hbf23de49,
32'hbefe3120,
32'h3d8ee592,
32'hbf784ff8,
32'h3c9173f6,
32'h3cd0c123,
32'hbea505ef,
32'h3dd8916c,
32'hbe8e1513,
32'hbe9f67a4,
32'hbf17bc94,
32'hbe10c274,
32'hbc256af4,
32'h3ed296b2,
32'h3e2f3c3c,
32'hbe0bccbc,
32'h3e94de47,
32'h3eb424dd,
32'hbdc6dd0c,
32'hbe06dd67,
32'hbe1223dc,
32'hbdcadbca,
32'hbc199fa2,
32'hbdeefba6,
32'hbd8cebcc,
32'hbbcc7d0f,
32'hbdecf6fe,
32'hbdd0fec0,
32'hbe58ad40,
32'hbdaa531b,
32'hbd8378c6,
32'h3a11f834,
32'hbd592ba0,
32'hbe9a0e5f,
32'hbe805520,
32'h3deba32b,
32'hbd7e4eb0,
32'h3e9b6435,
32'h3e36e16d,
32'hbf59f20f,
32'hbf23d87e,
32'h3c1cff64,
32'hbdd7d883,
32'h3e49ed81,
32'h3ede03d0,
32'hbe53de12,
32'h3e0db1f5,
32'h3e2187c4,
32'h3e348ece,
32'hbf04d1fa,
32'hbe645529,
32'hbd0b78eb,
32'hbd94b390,
32'h3e64470b,
32'hbd3d2728,
32'hbe2e8278,
32'hbebe267f,
32'hbbd57d13,
32'hbe42e610,
32'hbc4c790c,
32'hbda97652,
32'hbca09e74,
32'h3cf04fee,
32'hbf40769a,
32'hbf0b3442,
32'hbe23f478,
32'hbcb8481d,
32'h3de1eb12,
32'h3e90f8dd,
32'hbf81868a,
32'hbe843f19,
32'h3e673548,
32'hbeb4968f,
32'hbd5fa6e5,
32'h3dcfe8e0,
32'h3d4a8aa7,
32'h3d94a2d3,
32'h3e04af46,
32'hbdac3f72,
32'hbecc467d,
32'hbe021dd3,
32'hbd275e13,
32'h3c2f2bc5,
32'hbdd9b9c6,
32'hbe8019c2,
32'h3e02050c,
32'hbe5d9e06,
32'hbe5cd9ef,
32'hbda46525,
32'hbe206fbc,
32'h3ec5b957,
32'hbd0a6cac,
32'h3e62dc08,
32'hbf3fbcef,
32'hbee3a9fb,
32'hbd948ea3,
32'hbe08806d,
32'h3e8d0b7e,
32'h3e63e30f,
32'hbf713dfa,
32'hbe74f248,
32'hbd34049d,
32'h3cfbb00a,
32'hbcbd72b5,
32'h3c86f706,
32'h3e19fc99,
32'h3d58cd88,
32'h3d027dda,
32'hbc60bf0a,
32'hbee80c86,
32'h3df1ffa2,
32'hbc30b471,
32'h3cbbd604,
32'hbf0bff11,
32'hbee25baf,
32'h3dbacdf5,
32'h3d6e8872,
32'hbe3f55ca,
32'h3d2cbfc2,
32'hbe535dea,
32'h3c740ab5,
32'h3c177fdb,
32'h3cd858f6,
32'hbd4822d1,
32'hbdcfd972,
32'hbe294cd1,
32'hbe8263f8,
32'h3db1c01d,
32'h3d152b62,
32'hbefdcc7f,
32'hbee0efa9,
32'h3eb8cf46,
32'h3e61e246,
32'h3d936794,
32'h3d0c807e,
32'hbe3762bd,
32'hbe4fcdf1,
32'hbd8873c5,
32'hbdcf1c94,
32'hbeab3dc2,
32'h3d824ac6,
32'hbd4df357,
32'hbdbe6cd9,
32'hbf22a285,
32'hbed3aab6,
32'hbe2a8401,
32'h3d8a1780,
32'hbf08f654,
32'hbdb5525e,
32'hbe2560f4,
32'hbeeb41cd,
32'hbe693c81,
32'hbdf0afe9,
32'hbf251f32,
32'hbe1b9dc8,
32'hbc38ba38,
32'h3d8a820e,
32'h3e211059,
32'hbcf8e139,
32'hbf59222b,
32'hbedbdf7e,
32'h3d3b4208,
32'h3c3cf6e6,
32'h3dd97fae,
32'h3e8ff64e,
32'hbfcec6c8,
32'h3ceec108,
32'h3d5250c8,
32'hbe643a9d,
32'hbdce8c1c,
32'hbe3a72af,
32'h3d0e2d69,
32'hbcae3432,
32'hbeb074ee,
32'hbeaa3b38,
32'hbe89962e,
32'hbe5d029a,
32'hbe8fb55a,
32'h3d951e35,
32'hbe7d4096,
32'hbe88ac88,
32'hbe4f4a03,
32'hbdffdd32,
32'hbf4b675f,
32'hbd864fd4,
32'hbc729735,
32'hbe024895,
32'hbcdba17d,
32'h3d0565f5,
32'hbf947f39,
32'hbe99aa4b,
32'hbe1a6d91,
32'h3ea7da74,
32'h3d926ca6,
32'hbd917bfa,
32'hbf1d4cfa,
32'hbcf74b11,
32'h3e61de12,
32'h3e3a19ee,
32'hbe826002,
32'h3e71c12b,
32'hbdef5357,
32'hbd0f8872,
32'hbf03fedf,
32'hbeadda2e,
32'h3e4d8bc0,
32'h3e264747,
32'hbd47272b,
32'hbe6a7d41,
32'hbeebf773,
32'h3e934c55,
32'hbeb4aad3,
32'hbe06ab6b,
32'hbf1dc338,
32'h3b5b57fe,
32'hbe262503,
32'hbc02dd91,
32'h3e42b4ae,
32'h3d896f43,
32'hbf1b3ee2,
32'hbdbce0dd,
32'h3ede5407,
32'h3e82a475,
32'hbec58327,
32'hbdb0ef54,
32'hbfa991a1,
32'hbd93d391,
32'h3d88e29e,
32'hbd7a7090,
32'hbea29238,
32'h3e5d6de3,
32'hbd569ada,
32'hbde85e08,
32'hbfa9f73f,
32'hbf00ff6e,
32'h3c813c67,
32'hbaaacabd,
32'h3eaa0753,
32'h3d21ac40,
32'hbed44156,
32'hbe9f1b5b,
32'h3ec77fd0,
32'h3cc672ac,
32'hbf042fba,
32'hbe8a753b,
32'h3e2fe389,
32'hbe2ab24b,
32'h3d0e1142,
32'hbce60645,
32'hbf2398ea,
32'hbe25d47e,
32'hbeaf76df,
32'h3eff8451,
32'hbeb75c30,
32'hbb877950,
32'hbfe71063,
32'h3e7aa8d5,
32'hbed402dc,
32'hbe9faa1a,
32'hbefccbd2,
32'h3e17239f,
32'hbca9a567,
32'hbbcc0393,
32'hbf5ae729,
32'hbe0ae140,
32'h3eb82fee,
32'h3be1ebb5,
32'h3b8e9d5c,
32'hbe3f2a5e,
32'hbe882b03,
32'hbd6735aa,
32'h3e7eaf2b,
32'hbc9b573a,
32'hbf3ca028,
32'hbcf3ab8a,
32'hbe450827,
32'hbe851e6f,
32'h3da0017c,
32'hbecf9e6a,
32'hbf842a69,
32'hbc4fc3ca,
32'hbec559d1,
32'hbd3c5b0d,
32'h3ebab925,
32'hbe4c49f8,
32'hbf0bae2e,
32'h3e93c6d1,
32'hbe18b34b,
32'hbef9ece1,
32'hbe885cd9,
32'h3e767b56,
32'hbc819df0,
32'h3d784a69,
32'hbf4dc7e5,
32'hbeace7b7,
32'h3e868bf6,
32'h3c3a8be4,
32'h3e0b20cc,
32'h3da5780b,
32'hbe732156,
32'h3e9850a8,
32'h3ea78f36,
32'hbf074c2d,
32'hbec0daec,
32'hbe2c6dab,
32'hbcb2f9b7,
32'h3dab0a58,
32'hbe2dde60,
32'hbc889f39,
32'hbe907abe,
32'h3ed4d030,
32'h3d8b636e,
32'h3bc604e6,
32'h3e285036,
32'hbf7bdb59,
32'h3db33070,
32'h3bd3c40b,
32'h3e8a2048,
32'hbf3a1fa9,
32'hbfa4b4f0,
32'hbee71cfd,
32'h3ca5e8f9,
32'hbc99c49f,
32'hbf5dc1e9,
32'hbe5fd504,
32'h3ed69062,
32'h3dc4ff54,
32'h3e82743c,
32'hbe664080,
32'hbe57accf,
32'h3ea1c8e0,
32'hbe360751,
32'hbe864b9c,
32'hbd1646d5,
32'h3ba1d803,
32'hbcc2762b,
32'hbf8f1d10,
32'hbe03f667,
32'h3e6a99ee,
32'hbe340b2f,
32'hbdc8a47f,
32'hbefd107e,
32'h3e8876b6,
32'hbe76253a,
32'hbf5ca29a,
32'h3eb7743b,
32'h3ebd97b9,
32'h3db94022,
32'hbf949c65,
32'hbeeaad36,
32'h3ddf869e,
32'hb9b02880,
32'hbdcb3b34,
32'hbf6667a4,
32'h3e040080,
32'h3c19a770,
32'h3e1cf762,
32'h3d7a0f88,
32'hbe9bee40,
32'hbeb791dc,
32'hbdf2deb5,
32'hbed81f6b,
32'h3d268380,
32'hbe9a6b28,
32'hbeca5837,
32'hbccbb7ca,
32'hbf03a41a,
32'h3e8ab770,
32'h3e68dbc9,
32'hbf68a1f3,
32'h3f150f44,
32'hbe0dab76,
32'hbe05b59d,
32'hbd52526f,
32'hbf58d5ec,
32'h3dec4d20,
32'hbea511b4,
32'h3b7950e9,
32'hbfc72b30,
32'hbe4317a4,
32'hbf017341,
32'hbd10e105,
32'h3d8a60c9,
32'hbf564835,
32'h3edd3bfc,
32'h3e825587,
32'h3e280900,
32'h3e3e05cf,
32'h3e9eeeab,
32'hbd81a523,
32'h3e14f517,
32'hbe76696d,
32'hbdd83896,
32'hbc849344,
32'hbefb1445,
32'hbe8aac42,
32'hbef2edd7,
32'h3e2f65b4,
32'hbe07802c,
32'hbf36ca8c,
32'h3ee12e3c,
32'h3d939fee,
32'hbeb134d8,
32'h3d5df4ab,
32'hbef4df14,
32'h3d9b0b2f,
32'h3dfc8643,
32'hbea863c6,
32'hbf8b7be3,
32'hbf88548a,
32'hbd862690,
32'hbb009cc4,
32'hbcd5ba11,
32'hbf297c3d,
32'h3f4f2ce7,
32'h3ef33122,
32'h3e7c62dc,
32'h3f2b5243,
32'h3db086c9,
32'hbde12351,
32'hbf12f5ef,
32'h3f4f720c,
32'hbe05e692,
32'hbf6e6383,
32'hbebdb129,
32'h3e62c194,
32'h3e050dfe,
32'h3f45adde,
32'hbdb01816,
32'hbb25317b,
32'hbf0fef5a,
32'h3dceb7d0,
32'hbf900896,
32'h3f18710d,
32'hbfbffa84,
32'hbd6abee7,
32'hbe99df35,
32'hbe020616,
32'hbf1b789d,
32'hbef6d490,
32'hbe03caf6,
32'hbd9a9cc6,
32'h3d497b40,
32'hbf301676,
32'hbe0a21ed,
32'h3f1a182a,
32'h3e1127c5,
32'hbf1d9dde,
32'hbe60972e,
32'hbe425ad5,
32'h3d910ee6,
32'h3f5786d8,
32'h3e1b6a29,
32'hbf07119b,
32'h3d8c5426,
32'h3cfbdebf,
32'hbf3500ff,
32'h3ecefb4d,
32'h3d71deb7,
32'hbf2a8dd8,
32'hbf20ea1f,
32'h3f004c4c,
32'hbda82549,
32'h3f117cdb,
32'h3e86cabd,
32'h3f0a8bdc,
32'hbf901e82,
32'hbf28defe,
32'hbea9b3f5,
32'h3d2432c4,
32'hbe163d63,
32'hbc2fa703,
32'hbcb0d8a3,
32'hbee87c3e,
32'hbec46b43,
32'h3f02acc7,
32'h3f89a3a3,
32'h3fa6ef00,
32'hbeb06565,
32'hbf1c9424,
32'h3c1ef372,
32'h3e773f74,
32'hbb639949,
32'hbe072c71,
32'h3f3090b5,
32'hbf1e191c,
32'h3f966e5c,
32'h3eb97bb2,
32'hbd6e7a8f,
32'hbf3c91ef,
32'h3de24cb6,
32'h3ea5d9fa,
32'hbd9aac55,
32'h3d160051,
32'h3f249d8a,
32'h3dddc9ca,
32'hbef682b0,
32'hbf26198c,
32'hbe76da1e,
32'hbe283501,
32'h3dd6fe70,
32'h3bffb70b,
32'h3a325849,
32'h3f1c90c1,
32'hbfb25b40,
32'h3d2aaaa0,
32'h3f97b821,
32'h3f6702f9,
32'h3f4e8011,
32'h3ea609b0,
32'h3ec9c49e,
32'h3f7d14e4,
32'hbf1c5993,
32'hbda24d14,
32'h3f8b7a6d,
32'hbf105151,
32'h3f04a5b4,
32'hbe107634,
32'h3eb06692,
32'hbef02b91,
32'h3eea43d6,
32'h3f8a9734,
32'h3d1a052c,
32'hbea527d3,
32'h3efc75cd,
32'h3e2b50ad,
32'h3e8da1f3,
32'hbe11115c,
32'hbe58a63c,
32'hbe9ed76f,
32'h3f8a1525,
32'hbd3440d9,
32'h3d52be60,
32'h3f716812,
32'hbfc10704,
32'hbe6ca7e3,
32'h3e4bae87,
32'h3ed99423,
32'h3f59fba4,
32'hbeac6fbd,
32'h3f448d9f,
32'h3f1d3b2d,
32'hbf2411ce,
32'hbcd47047,
32'h3d50255c,
32'hbd49673a,
32'hbc5de722,
32'hbf31e51b,
32'h3ce141a1,
32'hbf308e4c,
32'h3f587f30,
32'hba9f7d2e,
32'h3d291ac4,
32'hbc95c2b7,
32'hbd8ac442,
32'h3d2739e1,
32'hbdb41a35,
32'hbd45617e,
32'h3d4fc70a,
32'hbd3fee90,
32'hbddd68eb,
32'h3d80296d,
32'h3dd0c93f,
32'h3d18a80d,
32'h3d8ffe8e,
32'h3cc44792,
32'hbce4eaaf,
32'h3d506388,
32'h3daab4db,
32'hbbdd00d4,
32'h3dbc948e,
32'h3c815dd4,
32'h3a387199,
32'hbceee2cd,
32'h3d830fbe,
32'h3d09eb11,
32'h3c68c6c5,
32'hbd847c1e,
32'hbbe280a1,
32'h3daddb18,
32'h3d8eff72,
32'h3d0ce43b,
32'h3d38a17b,
32'hbd808fd5,
32'h3c84aa69,
32'hbd89b832,
32'hbcd3452b,
32'h3dda342e,
32'hbd39ee17,
32'hbc8ea90d,
32'h3c51e3d9,
32'hbd63a0b9,
32'h3d81c4ba,
32'hb99779af,
32'h3d5630c4,
32'hbb965ac3,
32'hbc9f91f6,
32'hbd751b7e,
32'hbdc4cf28,
32'h3d95ef1f,
32'hbdae6333,
32'h3b1ec166,
32'hbd309c1a,
32'hbcb48f2f,
32'hbc880e84,
32'hbc534af1,
32'hbdb5bca0,
32'h3b8dc968,
32'hbb8b8a16,
32'hbd2029b5,
32'h3daa50e7,
32'h3cc36c75,
32'hbd1bdcdf,
32'hbcbd1cb2,
32'hbc9a1a3e,
32'h3cc559db,
32'hbb648ac2,
32'h3ca55ff5,
32'h3c59830e,
32'h3d9b9208,
32'h3d322204,
32'hbb5bffe2,
32'h3bbb99eb,
32'h3daa8b17,
32'h3cf76299,
32'h3de6dd2f,
32'h3d1ea977,
32'h3d4f2898,
32'hbc8c3f99,
32'h3dbfa969,
32'h3db32a98,
32'hbccfbae1,
32'hbc0a60c3,
32'h3dd9665e,
32'hbdc20530,
32'hba5b2a2a,
32'h3d68799e,
32'h3dde8580,
32'hbd266e21,
32'hbd08ff11,
32'hbd775d3a,
32'hbc167ac8,
32'h3da13fc3,
32'h3ec6a35b,
32'h3c0de8fa,
32'h3e46dbbe,
32'hbe9cf30d,
32'h3eb596e3,
32'h3db180c7,
32'h3c6928c7,
32'h3cb12fc2,
32'hbce7e1f4,
32'h3d464369,
32'h3d581e70,
32'h3e3a9893,
32'hbe0e2863,
32'hbe0106bc,
32'hbd6de5b8,
32'h3d353a17,
32'hbdadf984,
32'hbd7d6a04,
32'hbdf177c2,
32'hbe5e3af2,
32'hbd4c1fb1,
32'hbe90d146,
32'hbd3c1e9a,
32'hbdfd9884,
32'h3e548f77,
32'hbc90f513,
32'hbe3c6c64,
32'hbe76a69a,
32'hbef94b73,
32'hbe0e6839,
32'hbeb0fb95,
32'h3dcdceba,
32'hbec1464d,
32'hbe3114d7,
32'h3e9479b2,
32'hbeb137ed,
32'hbf24740d,
32'hbc5042d7,
32'hbc0f5056,
32'hbca123f2,
32'hbea5eaa8,
32'hbfabdf47,
32'hbdae8eee,
32'hbf89ae26,
32'hbe895317,
32'h3cbf3301,
32'hbf2ecd74,
32'hbcae8ad0,
32'hbe48c2d9,
32'h3ea189ab,
32'hbe43de23,
32'hbeda18cd,
32'h3f257234,
32'h3d3ce043,
32'h3f7c90f7,
32'h3c2103bd,
32'h3e6cadaa,
32'hbcdf7c7f,
32'hbe19acb4,
32'hbea58047,
32'hbed29a21,
32'h3ef7f54e,
32'h3eed8697,
32'h3f768d3a,
32'h3db9af98,
32'hbde7a5e0,
32'hbf465678,
32'h3d3de5f4,
32'hbb2237f7,
32'h3d7fccaa,
32'hbf70a38e,
32'hbf8d0f95,
32'h3e36ead6,
32'hbedfcb57,
32'hbf0bac7e,
32'hbec44efe,
32'hc00278ef,
32'hbea0f0c4,
32'hbef4d67d,
32'h3f1a1548,
32'hbcc60b9e,
32'hbf1058ba,
32'h3f554444,
32'h3f5ad0fb,
32'h3ed2375a,
32'hbe3ff92c,
32'hbd07fd6c,
32'h3d56a2ca,
32'h3eca7b6b,
32'h3e819657,
32'hbea47df5,
32'h3f68699c,
32'h3eb7bd58,
32'h3f4f3a3a,
32'hbdcaeb4a,
32'h3da0df2f,
32'hbf9344ea,
32'hbe9994a2,
32'h3dbcbeed,
32'hbdd1843f,
32'hbf70a671,
32'hbf789b7f,
32'h3e84a07a,
32'hbd03a3a0,
32'hbee204bb,
32'h3e4a4373,
32'hbf15ae47,
32'h3db7ed45,
32'hbec5cddd,
32'h3f1a444e,
32'hbd2be0b4,
32'hbf056628,
32'h3ec66cfe,
32'h3f691849,
32'h3ec48e59,
32'h3ed97c00,
32'hbf346bc7,
32'h3f02d781,
32'hbd3bc3b3,
32'h3e01be78,
32'hbe938cc4,
32'h3ef13f45,
32'h3f0bd16e,
32'h3d12a2ce,
32'h3e43ecdb,
32'hbe870886,
32'hbf1c71e2,
32'h3f55a1c7,
32'hbc3a2541,
32'h3d923539,
32'hbfafe7ee,
32'hbfc87bf8,
32'hbe2a564d,
32'hbc0c8fb7,
32'hbf4472b7,
32'h3f3ace22,
32'hbf77f847,
32'hbd3b7d20,
32'h3dcf7747,
32'h3eeb2e19,
32'h3dbebdb5,
32'h3ea48e59,
32'h3eab33e6,
32'hbd59293b,
32'h3ce1bf6d,
32'hbdc06833,
32'hbf57b942,
32'hbf364119,
32'hbf021e6d,
32'h3ed22bbb,
32'hbe58e199,
32'h3da57924,
32'h3f17eeaf,
32'hbdcebf44,
32'h3d222907,
32'h3d77d756,
32'hbefb827b,
32'hbf12552c,
32'h3d3c2be8,
32'hbc1fb80f,
32'hbfa6967f,
32'hbf54f886,
32'hbe107b26,
32'hbe601d49,
32'hbf3f4cf6,
32'h3ed21e17,
32'h3de3997e,
32'hbf6fff95,
32'hbee41339,
32'h3eef6628,
32'h3db2ccc0,
32'hbe241fd9,
32'h3e55c351,
32'hbe22eaab,
32'h3de56fd5,
32'hbe8d2d3e,
32'hbf48426c,
32'hbf0c6a48,
32'hbee75bf5,
32'h3e37be2e,
32'h3e4bd0c9,
32'h3b3b12ce,
32'h3f13da5b,
32'hbe6545ac,
32'h3e7bd859,
32'h3e8e87bf,
32'hbec6b0a5,
32'hbf999bdb,
32'h3bbcf370,
32'h3c14a85e,
32'hbf763439,
32'hbf88d838,
32'hbf2fa831,
32'hbdd645db,
32'hbf216338,
32'hbe89dee7,
32'hbd051915,
32'hbe53b518,
32'hbeeb85be,
32'h3e00f8a6,
32'hbe08d5c9,
32'hbd6e6787,
32'h3e26a79c,
32'h3ebff804,
32'h3e03bcd0,
32'hbebe891a,
32'hbf0aa5c2,
32'hbe05025b,
32'hbbca3a80,
32'hbe9586e2,
32'h3e3e9a8d,
32'h3b4d34bb,
32'hbcfd0efe,
32'h3ea6d68d,
32'h3def80bd,
32'hbf43cc63,
32'hbf7a9fd2,
32'hbe0e07db,
32'h3dbf9bd6,
32'hbd770b92,
32'hbf7e2f63,
32'hbf56fc15,
32'hbf087f96,
32'hbeea6ab8,
32'h3ebc5c95,
32'h3ec4e703,
32'hbec5cf70,
32'h3ea78bc9,
32'hbda4dcf0,
32'h3cd98fb9,
32'hbfa032c3,
32'hbe81e2bb,
32'hbd1974f7,
32'h3d97d4de,
32'h3e4d17aa,
32'h3e2acfac,
32'hbf1ae677,
32'hbed4eb4d,
32'hbdb13a72,
32'h3de58b37,
32'hbecf12f8,
32'h3e004bbc,
32'h3dcbbc42,
32'h3d3003d3,
32'h3efe9534,
32'hbf1ca29a,
32'hbf61c83b,
32'hbe71abed,
32'hbd00070b,
32'h3c14054e,
32'hbf7fdef2,
32'hbef4a7dd,
32'hbf055d97,
32'hbcdac641,
32'hbe93311b,
32'hbe023423,
32'hbdec6726,
32'h3d2502d8,
32'hbe2a99b7,
32'h3dd3da7d,
32'hbf98d4e7,
32'h3e06ec50,
32'h3cf27e33,
32'hbcad11a9,
32'h3d4e8a6c,
32'h3c006697,
32'hbf354458,
32'hbd5c6fae,
32'hbde297d3,
32'h3e5b248b,
32'hbd4e3cec,
32'hbe6b4523,
32'h3eef7a3b,
32'hbe615726,
32'h3e82dba3,
32'hbf1f822a,
32'hbed8f08e,
32'hbe55f43b,
32'h3c0854ae,
32'h3d5752ce,
32'hbf423bd2,
32'hbee931d7,
32'hbd654ad3,
32'hbd3a2152,
32'hbd2bdffd,
32'hbe437f4a,
32'hbe116bfc,
32'h3ebd3758,
32'hbc8efa16,
32'hbd86eb07,
32'hbfc14df1,
32'hbc8b9c10,
32'h3e405632,
32'h3f069608,
32'h3e1b2bff,
32'h3e7f68ae,
32'hbe023c5c,
32'hbd4a4d83,
32'h3eddaea4,
32'hbba576d8,
32'h3e0f36ec,
32'h3ead5bd3,
32'h3f386237,
32'hbd1c9fee,
32'hbe83ebae,
32'hbf3277de,
32'hbdef1f0e,
32'hbe926b84,
32'hbd3b2000,
32'h3c0030cd,
32'hbe90e9a7,
32'hbf43575a,
32'h3d3d6ef9,
32'hbe44a9f2,
32'h3e9284d0,
32'h3e012fbb,
32'hbe8e3691,
32'h3dd81221,
32'hbd6ee0b4,
32'hbe5f7177,
32'hbfbf10f2,
32'h3da6e19d,
32'hbe890f80,
32'h3e597576,
32'h3e59e356,
32'h3de163e1,
32'h3e0d0e56,
32'hbedeebdb,
32'h3e0ea592,
32'hbc8c9e87,
32'hbe5d6d22,
32'h3df42225,
32'hbec86522,
32'hbe475518,
32'h3e9a35bd,
32'hbf2668d6,
32'hbf23ae22,
32'hbf4c93e3,
32'h3ce27019,
32'hbdcf2b40,
32'hbe3c4e60,
32'hbf3f7d5b,
32'h3d246a40,
32'hbe24aa4b,
32'h3e0e8715,
32'h3eb2d46d,
32'hbeb7e3cf,
32'h3e2e243a,
32'hbbe1fc9a,
32'h3dd09a58,
32'hbf713e44,
32'hbcc9ba35,
32'h3dcf2fbe,
32'hbd5264dc,
32'h3e9063ab,
32'h3e24278e,
32'hbed42afa,
32'h3e9b57ea,
32'h3eae2f8c,
32'h3e478f5e,
32'h3e67c4f2,
32'h3cc8d976,
32'hbf8b982c,
32'hbe0a2107,
32'h3e6d19f6,
32'hbef7c801,
32'hbecc1ef5,
32'hbf413770,
32'hbcc1535d,
32'h3d73dd07,
32'hbf3b6028,
32'hbf3bd941,
32'hbe91affd,
32'hbd3ae793,
32'h3de2c406,
32'h3ead6007,
32'hbf01dc0a,
32'h3e2caf34,
32'hbcfcdf26,
32'h3e228005,
32'hbfe94f30,
32'h3d8cc942,
32'hbddeb21c,
32'hbd42b083,
32'h3e908014,
32'h3e2c080c,
32'hbf739e61,
32'h3da7c2fb,
32'h3fb12fc7,
32'hbe37174d,
32'h3e3d96e6,
32'h3d01908c,
32'hbfd40a08,
32'h3c7295c4,
32'h3e3f4e8d,
32'hbebcde82,
32'hbc71cd47,
32'hbe93a5cf,
32'hbd8cd86d,
32'hbd6c9783,
32'hbf9bc194,
32'hbf3a73ba,
32'hbc9256ec,
32'hbc62cff0,
32'h3d836be6,
32'hbea50e87,
32'hbe8a6a43,
32'h3d9bdf77,
32'hbec4cedd,
32'h3d871fb9,
32'hbfb448f9,
32'hbc42783c,
32'hbd6a424e,
32'hbde908fc,
32'h3de6c77c,
32'h3c8c64ff,
32'hbefd456e,
32'hbe8cf416,
32'hbe625d2e,
32'h3e0dea67,
32'hbdc9abff,
32'hbe5fd4a1,
32'hbfcdf6c8,
32'hbf0594f6,
32'h3ca0ad4e,
32'hbf67ce88,
32'h3e1ba67e,
32'h3e019b97,
32'h3cd2c168,
32'hbc7a3e63,
32'hbfff06de,
32'hbf341d5f,
32'hbf110111,
32'hbcd5afe1,
32'h3e4d4570,
32'h3ee251e4,
32'hbe5d9a46,
32'h3e1ae944,
32'hbdafaf88,
32'hbe30b40d,
32'hbdc7a7d2,
32'h3e3d8eb4,
32'hbe15bbde,
32'hbecf2c03,
32'h3e1b74d6,
32'hbe983180,
32'hbf14c955,
32'hbdc0aa1c,
32'hbf8e15c6,
32'h3e7c6c69,
32'hbed1b56c,
32'hbed7abcb,
32'hbfb06b35,
32'hbe6df559,
32'hbd91b3b8,
32'hbe2d9a81,
32'h3eb4a115,
32'h3e71c464,
32'hbc56d157,
32'h3d2f0477,
32'hbff2c84e,
32'hbe71ec33,
32'hbd6ad431,
32'hbe9e6828,
32'h3e073359,
32'h3e1243aa,
32'hbe034b94,
32'hbdf0a3ca,
32'hbec410ca,
32'h3d684dea,
32'hbfe27e4a,
32'h3daf9912,
32'h3e87f448,
32'hbecbfd60,
32'h3e914804,
32'hbd8dd2b3,
32'hbee6b97f,
32'hbf084955,
32'hbfb327d3,
32'hbe8b8ea3,
32'hbaae5c16,
32'hbf807b1c,
32'hbfd185c8,
32'hbe727813,
32'hbe9de172,
32'hbe708926,
32'h3dd6beca,
32'hbf1958de,
32'hbd8e5848,
32'h3d2dff0f,
32'hc00ecfda,
32'hbee5d5ea,
32'hbe26acc0,
32'h38d5d1f5,
32'h3ed0ef31,
32'h3e9f3322,
32'hbdff14a6,
32'hbf1ef187,
32'h3cbea0ab,
32'h3e89c899,
32'hbfa3c723,
32'h3d2f4d3c,
32'hbf2f02c6,
32'hbf4325c3,
32'h3e4b932c,
32'h3e0631d4,
32'hbeb20ded,
32'h3f0cedbf,
32'hbfac7641,
32'hbe037fd2,
32'hbe4dcbae,
32'hbfa640e3,
32'hbf813e5c,
32'hbe00cd8a,
32'hbe3da659,
32'hbf9b7bbe,
32'hbf44f8ad,
32'hbf17f4de,
32'h3d70af94,
32'hbd1670c9,
32'hbff356d0,
32'hbf1cf13e,
32'h3f05b9d6,
32'h3e289e8e,
32'h3e5edd37,
32'hbe72597a,
32'hbc857852,
32'hbee493c5,
32'hbd80ede5,
32'h3e849ebd,
32'hbf92b234,
32'h3be4200b,
32'hbf18eb18,
32'hbf5fbd18,
32'h3da81707,
32'h3dcfd55e,
32'hbec2203c,
32'h3eb11ec9,
32'hbf8532e5,
32'h3e7bcb40,
32'hbe331d07,
32'hbfbceabe,
32'hbe6706a9,
32'hbf77c212,
32'hbda4a43b,
32'hbf60e32f,
32'hbe9bbe69,
32'hbf2b750d,
32'hbc763626,
32'hbc48982e,
32'hc000d23a,
32'hbebb0ede,
32'h3e53f2ba,
32'hbc22b865,
32'h3e8f989d,
32'h3dafbd28,
32'h3e45a151,
32'hbde21aaa,
32'h3e4afb0d,
32'h3e04681f,
32'hbf407a7a,
32'hbeca5171,
32'h3e547f57,
32'hbdcd72ce,
32'h3dfed233,
32'h3ed0de96,
32'hbef3bb86,
32'h3dbf61fd,
32'hbe85f68d,
32'h3b810082,
32'h3f71239d,
32'hbfb0be59,
32'hbdb10320,
32'hbfcbf6e9,
32'h3de291a0,
32'hbd141497,
32'hbe8a89a8,
32'hbf903fdf,
32'h3d343164,
32'hbc6ceef6,
32'hc0122daf,
32'hbe69611c,
32'h3fa19e0f,
32'h3ec7c507,
32'h3f5e6774,
32'h3ed3572f,
32'hbe358657,
32'hbebe2ab4,
32'h3f78f019,
32'h3ea785c9,
32'hbec18dd5,
32'hbe238ed0,
32'hbf37bd17,
32'hbfa370c8,
32'hbdbc72a1,
32'h3ec5bebf,
32'h3dd8743a,
32'hbdbce314,
32'h3e9f7568,
32'h3d3b8b8f,
32'h3f90c19d,
32'hbf95e9cc,
32'h3e4c443d,
32'hbe80d3ea,
32'h3f2f5718,
32'hbcce5f04,
32'h3da978a5,
32'hbf1acdaf,
32'hbd465bf1,
32'h3ce4342f,
32'hbf11d809,
32'h3e9e0fcb,
32'h3f118410,
32'hbe1c1bc4,
32'h3f18c496,
32'hbe35c6c9,
32'hbd46543f,
32'hbea62b83,
32'h3f423e7d,
32'h3f005ccd,
32'hbecbd441,
32'hbe2fbca3,
32'hbea99652,
32'h3de464df,
32'h3e90690f,
32'h3f342ff2,
32'h3e55b52a,
32'hbf2b83af,
32'h3f135816,
32'hbfa5d7e3,
32'h3f01337a,
32'hbfcd9403,
32'h3efa98b2,
32'hbf1757b1,
32'hbf1ac88f,
32'hbee99481,
32'h3db31273,
32'h3f2005c5,
32'h3ac3d500,
32'hbc82fc49,
32'hbf5d0fdf,
32'hbfc9aa40,
32'h3f0de197,
32'h3e940f65,
32'h3f6847a5,
32'hbe9c8e67,
32'h3f2ad3fa,
32'h3e5fa158,
32'h3ee6ebdd,
32'h3e22e76c,
32'hbef6faab,
32'hbefb2446,
32'hbcfc83f4,
32'hbedbec97,
32'hbd3fec0b,
32'hbd1ae832,
32'hbeb64174,
32'hbf016b3b,
32'h3ef6b9b5,
32'h3de99bed,
32'h3faed4aa,
32'hbe0e7005,
32'h3f00b54b,
32'hbf08b5b3,
32'h3cb18b04,
32'hbeb4f1bb,
32'h3f403d58,
32'h3ed5b8fb,
32'hbd99a514,
32'h3b99740f,
32'hbeb09f07,
32'h3f8b0086,
32'h3fba0e4a,
32'hbf23e7a0,
32'h400e6e09,
32'hbf8b549e,
32'hbfa39ca6,
32'hbf64c9f4,
32'hbf22386f,
32'h3eb523b3,
32'hbcc41ec8,
32'hbeb6a106,
32'h3fa08a51,
32'h3f21da02,
32'h3f6f2f5b,
32'hbf17ec9a,
32'hbd0313e1,
32'hbe9b6128,
32'hbd3982db,
32'h3b658ba2,
32'h3f7e01b2,
32'hbe1f9869,
32'h3f602472,
32'h3e8c2e48,
32'h3e1a43eb,
32'hbd9db51d,
32'h3eaf1ba4,
32'h3e966d92,
32'h3c81bc54,
32'h3dab5964,
32'hbf1bf8e1,
32'h3f5ac266,
32'h3f22a7c0,
32'h3e8f0001,
32'h3c2bf94b,
32'h3e2dd71a,
32'hbe7578f0,
32'hbddc217b,
32'h3f7c180b,
32'hbf34fb2e,
32'h3c9ff29b,
32'hbf1861d9,
32'h3f5c0ed0,
32'h3f0a3e14,
32'hbe82ca4b,
32'h3d4bae32,
32'h3d0bc5d8,
32'h3d89cbaa,
32'hbdd95c02,
32'h3db8e88a,
32'h3f3dd4ba,
32'hbbe8ba00,
32'hbd96314c,
32'h3e41ce17,
32'h3d254d02,
32'hbc0772d1,
32'h3d032d97,
32'h3e9b952b,
32'hbca714ff,
32'h3d372778,
32'hbcdaa203,
32'h3f5819e6,
32'h3ef044fe,
32'h3e8caf16,
32'h3d95442a,
32'hbbea792f,
32'hbe95bc30,
32'hbcbe3148,
32'hbdf1463c,
32'hbf01490e,
32'hbcc627ef,
32'hbf698331,
32'h3f639a64,
32'h3cd90498,
32'h3f215cc3,
32'hbe84c375,
32'h3b753052,
32'hbd35ca4a,
32'h3ddf30b4,
32'hbd945680,
32'hbd20c924,
32'hbc10eff6,
32'h3d5cb4a1,
32'hbcff58d8,
32'h384f00e9,
32'hbb50084b,
32'h3cbef4d1,
32'hbd8545df,
32'h3ce2b0da,
32'hbc1fd474,
32'hbd62dafd,
32'hbda044ca,
32'hbd34a3b7,
32'h3c3ec657,
32'hbce87816,
32'h3c9a34c5,
32'h3b1e14d5,
32'h3be035c7,
32'h3db5d201,
32'h3d66911b,
32'h3c868d45,
32'h3d81f072,
32'hbbea8723,
32'h3b114ddc,
32'hbc6cc889,
32'h3d6d4964,
32'hbbdd682f,
32'h3d919c83,
32'h3ca362d1,
32'h3baab996,
32'hbc7ddf6d,
32'h3d1fa428,
32'h3c80cff8,
32'h3d2dd121,
32'h3ccd4fe8,
32'h3c755c33,
32'hbc5158a4,
32'h3c0efd12,
32'h3ccdd567,
32'hbcc9dbb5,
32'hbd6ce35c,
32'h3d9d5cc4,
32'h3bd71687,
32'hbca67c58,
32'hbd6fd832,
32'h3c73600f,
32'h3d247bff,
32'hbcee8503,
32'hbdc03513,
32'hbbeba93d,
32'hbcf7a08d,
32'h3d392cc4,
32'hbd83036d,
32'hbb916540,
32'h3d0daaa1,
32'hbd38f52d,
32'h3dac6470,
32'hbcb069e2,
32'h3d2dec08,
32'h3c91aa35,
32'h3b0e47cf,
32'hbc2a2151,
32'hbb7ea99b,
32'h3cf16379,
32'h3d19afe2,
32'hbbe9f03b,
32'hbc4c2564,
32'hbc385df8,
32'hba092ce6,
32'hbd8731da,
32'h3d8f95cc,
32'h3d78090c,
32'h3cc1470f,
32'h3d928d02,
32'hbd4d35bd,
32'h3d8026ba,
32'hbd00281a,
32'hbcf8551f,
32'hbc31625f,
32'h3d3cf997,
32'h3dae89e8,
32'h3dc54422,
32'h3da941b4,
32'h3d0a1420,
32'hbcb0bb93,
32'hbd99154a,
32'hbcc4d46c,
32'h3baa148a,
32'hbcdc78e7,
32'h3e1b0195,
32'hbd56dd01,
32'hbd6ee40e,
32'hbcf41605,
32'hbe12e45a,
32'h3ea63a69,
32'hbd12184a,
32'hbcab3023,
32'h3d64e10d,
32'h3cc50f97,
32'h3cad5ff4,
32'hbd996c16,
32'h3dd8e604,
32'hbdd8e1f8,
32'h3bd8ec41,
32'hbda6019b,
32'h3d48dec1,
32'h3f13ef00,
32'hbebad3da,
32'h3b86aa72,
32'h3e171a82,
32'h3cea3088,
32'hbf4f833e,
32'h3e95132e,
32'hbdde5f9c,
32'h3ec8ff7c,
32'h3d64b347,
32'hbca900ce,
32'hbcaadb2c,
32'h3dfa9c7e,
32'hbc80dd36,
32'h3df43d08,
32'h3d500de7,
32'h3f937db1,
32'h3ebfac85,
32'h3c031abe,
32'hbe9f9860,
32'hbe2ff308,
32'hbcb49dc3,
32'hbc9813e0,
32'hbbfc9c41,
32'h3c15ceab,
32'hbddba05f,
32'h3ca96f63,
32'hbe9fd89b,
32'hbe49952b,
32'hbcb395bf,
32'h3e645e00,
32'h3d47d123,
32'hbd0f6770,
32'hbed87f39,
32'h3dd7ae0f,
32'hbd7fa677,
32'hbddbd0b5,
32'h3f426f5b,
32'hbf314bc6,
32'h3e03f3fb,
32'hbd1c6a9f,
32'hbe0bb568,
32'hbf194a7c,
32'h3f6fa6e0,
32'hbee625ef,
32'hbe9f01c9,
32'h3f7154d9,
32'h3d81518a,
32'h3fdb690f,
32'hbe988bde,
32'hbd49c528,
32'h3c45b1ef,
32'hb985aa93,
32'h3acc4604,
32'hbe53e12e,
32'hbe50c3f4,
32'hbec9484d,
32'h3f1ce9fd,
32'hbf5e421c,
32'hbed2db9d,
32'hbef1093a,
32'h3b36f8c3,
32'hbf366225,
32'h3eef88c8,
32'h3d145e26,
32'h3e218431,
32'h3f0297f9,
32'hbda4d108,
32'hbea45ece,
32'hbe123fdc,
32'hbde78868,
32'h3e266d28,
32'hbe81d765,
32'h3e9247ad,
32'hbf7f9539,
32'hbdec9d77,
32'h3f3eeb07,
32'hbe564bd7,
32'h3f3e75f3,
32'hbe5332b5,
32'hbe231709,
32'hbe0ddd69,
32'h3dbd0cda,
32'hbdb0d4fb,
32'hbfac18ac,
32'hbf941add,
32'hbe5b7f63,
32'hbe6a54bd,
32'hbf9db402,
32'hbf3e87ec,
32'hbe96d47b,
32'h3d8cdf3b,
32'hbf7222ba,
32'h3f096e30,
32'hbc933a4a,
32'h3f14377e,
32'h3e575548,
32'hbf7afc14,
32'h3e0210cf,
32'hbe122875,
32'hbe829bab,
32'h3e09ff04,
32'hbe97be1f,
32'h3eb8aa19,
32'hbe434060,
32'hbed8afaa,
32'h3e02a9f7,
32'hbe953588,
32'h3edba8bb,
32'h3d12a839,
32'hbf4241d9,
32'hbe404233,
32'h3d6fded4,
32'hbd20ef0f,
32'hbfc1dde9,
32'hbf5f61c1,
32'h3efefd0b,
32'hbf02de67,
32'hbfacdabc,
32'hbf0a98f7,
32'hbf482d65,
32'h3e707772,
32'hbf43b326,
32'h3f0b619a,
32'hbd0971db,
32'h3f72c8b9,
32'h3ed56688,
32'hbeac201a,
32'h3f2ace68,
32'h3d8953f4,
32'hbe992881,
32'h3dcc7548,
32'hbce8c162,
32'h3e85fbae,
32'hbcae01ca,
32'hbe658193,
32'h3eeca8f0,
32'hbf24b3e4,
32'h3f20981f,
32'h3e6f1be2,
32'hbf13389c,
32'hbeac5cbe,
32'hbd1921f4,
32'hbd8a40b8,
32'hbee6c305,
32'hbf6a9a27,
32'h3f427bde,
32'hbedf0c8e,
32'hbf8285d0,
32'hbf1473d4,
32'hbeb71937,
32'h3f361426,
32'hbf104655,
32'h3f6c3897,
32'h3c04a5a9,
32'h3f1d2722,
32'h3e981453,
32'h3e4a8056,
32'h3f1f64d1,
32'hbceaae4a,
32'hbee4e20d,
32'hbf6181c2,
32'h3f03244c,
32'h3e0958df,
32'h3eea0393,
32'hbf54a40b,
32'h3f0c9682,
32'hbeaa3273,
32'h3f4109df,
32'hbf5a3f19,
32'hbf098d84,
32'hbde8035c,
32'hbd97d008,
32'hbc01cc32,
32'hbcae9512,
32'hbfac54b7,
32'h3f1af9ea,
32'h3dad23b1,
32'hbe71ecbe,
32'hbed0d7ae,
32'hbd96d6df,
32'h3e2d58de,
32'hbec98225,
32'h3f0746b0,
32'hbcbcc13d,
32'h3d7b1188,
32'h3ef80344,
32'h3eac3037,
32'h3ef4ac77,
32'hbebd3b40,
32'hbf35f8e6,
32'hbf39152e,
32'h3e5c7cf1,
32'h3e92045a,
32'h3e025c44,
32'hbf83fd71,
32'h3d51081c,
32'h3de9c08a,
32'hbeb4d92e,
32'hbfd99396,
32'hbfc05053,
32'hbe0abaa3,
32'h3d7d5ac8,
32'hbc7144ac,
32'hbfe79af7,
32'hbfaec2ab,
32'hbeb558c0,
32'hbe22c984,
32'hbe0ed296,
32'hbecf0456,
32'h3db40fcb,
32'hbf93781f,
32'hbdbd25bb,
32'h3f3223f0,
32'hbd1ab9d0,
32'h3e60f4af,
32'h3e111cfa,
32'h3e7bab1c,
32'h3ef5e529,
32'hbde63c59,
32'hbf192a8c,
32'hbf787246,
32'hbcb65291,
32'h3e82d3cf,
32'hbd076222,
32'hbf9aad12,
32'h3d6adf9a,
32'h3e3363d8,
32'h3efd9f23,
32'hbf0e59b5,
32'hbf789515,
32'hc00da2ba,
32'h3d8f2a92,
32'h3cc25aee,
32'hbf84453c,
32'hbfa2a1f7,
32'hbf7773ec,
32'hbe4082c2,
32'hbf774a9a,
32'hbe7132d6,
32'hbec7541b,
32'hbeacfdc1,
32'hbe2b33e2,
32'h3ef2db30,
32'h3bff9bcc,
32'h3ec47da9,
32'h3e6dcd38,
32'hbe0ceb92,
32'h3ec06a3d,
32'h3e7ee1ea,
32'hbe988b40,
32'hbf523800,
32'h3e9413bc,
32'h3e9af6a1,
32'h3de00cd8,
32'hbfafae37,
32'h3ece8387,
32'h3dd2c83a,
32'h3dcb1553,
32'h3daaa721,
32'h3ebcaa5c,
32'hbff6da39,
32'h3d8b6ff5,
32'h3d102520,
32'hbfb27586,
32'hbf7dd6c3,
32'hbeff0e09,
32'hbeaa3b6f,
32'hbf7cb63a,
32'h3d235b76,
32'hbe38abff,
32'hbea918b2,
32'hbec09ccf,
32'h3e8adc07,
32'h3e803700,
32'h3e20bb5b,
32'hbd4c3622,
32'h3cc77128,
32'h3ea04ed4,
32'h3c97625a,
32'h3d0601c9,
32'hbf41faf4,
32'h3e3e58a3,
32'h3e7b69f1,
32'h3ee92ec2,
32'hbf62cfe6,
32'h3e0a8c42,
32'h3f1e6abc,
32'hbe729f17,
32'h3d7cb946,
32'h3e8b37c2,
32'hbfe8d802,
32'hbdb1a30d,
32'h3c8444fc,
32'hc0072126,
32'hbf5aed2b,
32'h3ee6cb93,
32'hbeb66e0e,
32'hbfa85b55,
32'hbce05124,
32'hbca888ad,
32'hbe934493,
32'hbe8eb051,
32'h3e1b93b8,
32'hbe2bcd10,
32'hbe9ec7ed,
32'h3e4e0df7,
32'h3e98633a,
32'h3e9bb89b,
32'h3b2d14e1,
32'hbed47eb1,
32'hbfc80221,
32'h3dc48bc9,
32'h3c40721d,
32'hbdb13535,
32'hbfac862b,
32'hbf56acce,
32'hbeb4b002,
32'h3f06630a,
32'hbe1c5307,
32'hbe8cd2a1,
32'hbf5e0147,
32'h3d7ee954,
32'h3cca560c,
32'hc0010b8c,
32'hbf72bf3c,
32'h3eae72a1,
32'hbd01c4c4,
32'hbee45bcc,
32'hbed8209f,
32'h3d2c715c,
32'hbe634b4d,
32'hbd9829e5,
32'h3e8ca50e,
32'hbf097b5f,
32'hbe8e43c8,
32'hbe26531a,
32'h3d6da1fd,
32'h3ede6b97,
32'h3d95cf16,
32'hbf1de47c,
32'hbeff63d7,
32'h3eb32d76,
32'h3ecae50d,
32'h3e65a70c,
32'hbfc21999,
32'hbfd6fd8e,
32'hbea037e9,
32'h3e9186df,
32'h3e8bee6f,
32'h3c5b428f,
32'h3e9013a4,
32'h3d8b5b12,
32'hbd75e76c,
32'hbfeb588b,
32'hbf84e5c9,
32'h3e667658,
32'h3d047b5c,
32'h3e18eb86,
32'hbe137073,
32'h3dd3ca80,
32'hbeb4a187,
32'hbd4f7330,
32'hbc0a9241,
32'hbf337791,
32'hbe1853f6,
32'hbec85cc8,
32'h3df61d0a,
32'h3e439fec,
32'h3d929a56,
32'hbe90c38c,
32'hbf53beaa,
32'h3c2a585b,
32'hbe1a776a,
32'h3ed58945,
32'hbf75e037,
32'hbff9f36d,
32'hbde82108,
32'hbea92c89,
32'h3eaa0e81,
32'hbdb27081,
32'hbf72602a,
32'h3d558511,
32'h3caed09c,
32'hbfc67c46,
32'hbffe0ab9,
32'hbf398235,
32'hbe9e690d,
32'h3f369b92,
32'hbe00a4f7,
32'hbd434c91,
32'h3e7d66c6,
32'h3c9ca323,
32'h3e5f26f4,
32'hbe88d5c6,
32'h3ef65da7,
32'hbea0db5b,
32'h3e97d67d,
32'h3edc5cc3,
32'hbd546e6b,
32'h3eb4f68e,
32'hbf31d4fd,
32'hbf6a1d8e,
32'h3e9d18ea,
32'h3e846445,
32'hc023e397,
32'hbfd043e0,
32'hbf07ddc8,
32'h3e87368a,
32'h3cd12743,
32'h3e94594f,
32'hbfdb0055,
32'hbcfec3f2,
32'hbda75260,
32'hbfa07711,
32'hbf67b591,
32'h3e3017bd,
32'hbe2df59b,
32'hbf0821b6,
32'hbee3021d,
32'h3bbcbcc7,
32'hbe8c037a,
32'hbef69534,
32'h3ea777a3,
32'hbf517278,
32'h3e99057c,
32'hbe1d23eb,
32'h3ee066bb,
32'h3eca0411,
32'hbe8056fe,
32'h3e7a5aed,
32'hbf9efac6,
32'hbf1d9039,
32'h3e8b42d0,
32'hbe2ef522,
32'hc030d317,
32'hbed4aa3e,
32'hbeb941eb,
32'h3e570c43,
32'h3dd292cd,
32'h3e14721b,
32'hbf83b624,
32'hba0b6600,
32'hbd2bee81,
32'hc01371ba,
32'hbebf2f21,
32'hbe9fa3ff,
32'hba501356,
32'hbf1c3f89,
32'h3e8b2d00,
32'hbe5c6ca5,
32'hbea4b6f4,
32'hbebe8aee,
32'h3f63675a,
32'hbdecbe49,
32'h3d88451a,
32'hbe8f5dcb,
32'h3bbcbebb,
32'h3e8df759,
32'h3f3d5685,
32'h3f127284,
32'hbf7eb247,
32'hbf356c91,
32'hbe8aca12,
32'hbee10498,
32'hc0299ad2,
32'h3e19211a,
32'hbf6ac04a,
32'h3eb2ba6d,
32'h3e6a3a3e,
32'hbed1979a,
32'hbf44e646,
32'h3b1918d1,
32'h3d8ffeb0,
32'hbffdf40f,
32'h3ec35913,
32'hbe6755cf,
32'h3ea2e0c4,
32'hbf016787,
32'h3e650e71,
32'h3e50f771,
32'hbf303a1a,
32'hbd6e0dc3,
32'h3e95c0e6,
32'hbd07e8c7,
32'hbdf9183d,
32'h3dc906d0,
32'h3e971bde,
32'h3e016fc2,
32'h3f1f445b,
32'h3f0e2d82,
32'hbee29437,
32'hbeec7848,
32'h3f2295aa,
32'hbe88aca6,
32'hc02d1878,
32'hbec0aa46,
32'hbf3ad8e5,
32'h4008ce64,
32'h3ef6efad,
32'hbe52c25d,
32'hbee656c0,
32'h3c97a888,
32'hbc0e60ea,
32'hbfefa502,
32'hbec0945c,
32'hbe67214d,
32'hbecf42a5,
32'hbeef0144,
32'hbedc1ca7,
32'hbe9d18b4,
32'hbec7a153,
32'hbf0ab76c,
32'h3e6f9df9,
32'hbf55bf3b,
32'h3eb62416,
32'h3e835fff,
32'hbea8a5a0,
32'h3f437fda,
32'h3ebd9b96,
32'hbe01dcab,
32'hbfd544d5,
32'hbe1c7546,
32'h3eba4df7,
32'hbe9b502e,
32'hbfb886bc,
32'h3eb80a00,
32'h3e4256ee,
32'h3e1a08dc,
32'h3f374716,
32'hbe17b5d9,
32'hbed65c5e,
32'hbca50cd2,
32'hbb89b9e8,
32'hbf9ff2b6,
32'hbf84c6f1,
32'h3ed3972a,
32'hbe09d4e5,
32'h3f48b3e3,
32'hbeed0e39,
32'h3c293177,
32'hbf20737d,
32'h3edf976d,
32'hbe081091,
32'hbdf7cca9,
32'h3eb6f074,
32'h3ea57ce4,
32'hbf85ee24,
32'h3d1fe944,
32'hbe524d07,
32'hbe7834ea,
32'hbfb602c7,
32'hbe41108e,
32'h3f404742,
32'hbee658ad,
32'hbf658380,
32'hbe499945,
32'hbdd4b401,
32'hbedb8be4,
32'h3f213078,
32'hbebc6f9d,
32'h3d9d08ec,
32'hbcf2c644,
32'hbdb59a44,
32'hbfc0e6de,
32'hbf842220,
32'hbd6af31d,
32'hbf084e77,
32'hbe86d2a7,
32'hbf243d79,
32'hbea2bb7b,
32'hbef59084,
32'h3df1216c,
32'h3ee14fee,
32'hbcd10b5c,
32'h3f06885a,
32'hbf0ffc14,
32'hbf947612,
32'h3d1ba11d,
32'h3e98556f,
32'hbee100af,
32'hbfcc6d22,
32'h3ecf0d1e,
32'h3dabc70f,
32'hbfa0f7b1,
32'hbf7b6849,
32'h3d5b8c48,
32'hbe2138bf,
32'hbf1fec49,
32'h3f22fa23,
32'hbee9ba15,
32'h3e27339a,
32'hbd0eb3fa,
32'h3a861cf4,
32'hbf562165,
32'hbf268d17,
32'hbd9fcf40,
32'hbf8abd28,
32'hbe1a014d,
32'hbe6bdebf,
32'hbf8a019d,
32'hbf819fa5,
32'h3ec05931,
32'h3f7e2bf3,
32'hbd642556,
32'h3f3902c7,
32'hbf6d06e2,
32'hbf30b481,
32'h3e2bf09d,
32'h3ef1b310,
32'hbe5bc09a,
32'hbefcda1c,
32'hbf988f12,
32'hbebdcba3,
32'hbf8b247f,
32'hbf9de506,
32'h3ceb0281,
32'hbf0b43aa,
32'hbf87f608,
32'hbf91a9a2,
32'hbe71df6c,
32'hbd807e7b,
32'hbd3de63b,
32'h3b73d4c5,
32'h3f014464,
32'hbe053eb8,
32'h3e71d77d,
32'hbf8b9a74,
32'hbe463c69,
32'h3eca94f9,
32'hbe2ac428,
32'hbe8ee758,
32'h3f8f663b,
32'h3f149b97,
32'hbd647dd6,
32'h3db5acb6,
32'h3e94fc02,
32'hbea8aaf2,
32'hbf815634,
32'hbd972da8,
32'hbd9fb4f4,
32'h3e4e5825,
32'hbdb38b16,
32'h3d3031ab,
32'hbf095380,
32'hbec0f227,
32'hbebb5730,
32'hbcd46e81,
32'hbc33fe8f,
32'h3d07e7cf,
32'h3d7a9905,
32'hbddbcdac,
32'hbd279a48,
32'hbd34cbcd,
32'h3e12a0a7,
32'h3f3b869a,
32'h3f052694,
32'hbfc69b81,
32'hbc6542d3,
32'hbe8ddf78,
32'hbef1c108,
32'hbf3b89e0,
32'hbe9ab116,
32'h3fbca837,
32'h3c826799,
32'hbe3d3be4,
32'h3ed01d5f,
32'h3ee4e7a7,
32'h3eaf1205,
32'hbe2056d1,
32'hbd7af515,
32'hbf3a6748,
32'hbd154714,
32'hbc944c02,
32'h3e9ed049,
32'hbd9ca709,
32'hbb7e1057,
32'hbd618c43,
32'hbdb0d2a7,
32'h3d53e21e,
32'h3dc0d87e,
32'hbd32ab10,
32'hbd22563e,
32'hbd87a0f1,
32'hbd5931a9,
32'h3f485635,
32'h3ef41ee1,
32'h3e324d1a,
32'hbc893770,
32'hbdc377aa,
32'h3f098107,
32'hbdc5a2b9,
32'hbd99699a,
32'hbf5caf5c,
32'hbcb986bb,
32'hbea01876,
32'h3f0bc359,
32'hbdb8ee6e,
32'hbe32d889,
32'hbd6fd9dd,
32'h3adadf76,
32'hbd9015f2,
32'h3d2a1baa,
32'h3de40d71,
32'h3f3d923e,
32'h3d8c6a3d,
32'h3ce56783,
32'h39dc0282,
32'h3d9e859b,
32'hbc870b8b,
32'h3da18b7a,
32'hbd505769,
32'h3d0c4388,
32'h3d7f0c1c,
32'h3d2d53e1,
32'h3f5c7457,
32'h3f1cc154,
32'h3e85c4cb,
32'h3d835560,
32'h3c944f0c,
32'hbeaf7c88,
32'h3b8323a9,
32'hbd7a75bb,
32'hbe89d04b,
32'h3c51aa9a,
32'hbf50c76d,
32'h3f42c41d,
32'h3d8ac586,
32'h3f2f5719,
32'h3d5f865e,
32'hbd73a8e3,
32'hbdb8966b,
32'hbd81ae7a,
32'hbd888d49,
32'h3dbfdbbc,
32'h3d266db0,
32'hbca0fe22,
32'hbaa462ae,
32'hbd2d87b6,
32'hbc06c34a,
32'h3d8f684f,
32'hbcd8cca3,
32'hba6db97d,
32'hbd13f4ea,
32'h3bb75046,
32'h3db74af6,
32'hbd3f3854,
32'hbbe80fd7,
32'h3d33d8e7,
32'h3d74da88,
32'hbd460f5c,
32'hbcb7d226,
32'hbb1985f0,
32'h3d3c54bd,
32'hbd98f8b0,
32'hbbe01604,
32'h3ca6a36e,
32'hbd6501fd,
32'hbde16b65,
32'h3cbea478,
32'h3b882000,
32'hbd6f0ac0,
32'hbda1a6f9,
32'h3d6767e2,
32'h3d9ac9db,
32'hbc1af644,
32'hbdaf2d57,
32'hbdab6435,
32'h3d788eab,
32'h3db61100,
32'hbda337a1,
32'h3d3b6ae3,
32'hbd4702ec,
32'h3c247aa9,
32'hbd2212c0,
32'h3d4757f6,
32'h3d7dbc1d,
32'h3dd544ee,
32'hbc2d6593,
32'hbdc43455,
32'h3ddc9dd7,
32'hbd46ca92,
32'hbc84a6a9,
32'h3d89ddf2,
32'hbd22a905,
32'hbcab70ea,
32'hbc05e09f,
32'hbc85d592,
32'hbd36bd71,
32'h3d82d3ba,
32'h3d1b7976,
32'h3b0b58ac,
32'h3c8f1c36,
32'h3c6dd145,
32'hbd738837,
32'h3aab4c5f,
32'h3d754b2b,
32'h3cb9ae99,
32'h3d0d537f,
32'hbc825b7f,
32'hbd18d327,
32'h3da626d3,
32'hbc900068,
32'h3d0bb5e6,
32'h3c63ab52,
32'hbc8ed068,
32'h3cbef4a5,
32'h3dbae513,
32'h3adf687f,
32'hbc55dffd,
32'hbc933608,
32'h3d901563,
32'hbc7013dd,
32'h3d35ec41,
32'hbd81aa01,
32'h3d8d00bd,
32'hbd7a5f91,
32'h3d9b5408,
32'hbc5ac818,
32'h3d76ebac,
32'hbd0c95ac,
32'hbd4351b2,
32'h3d302d96,
32'h3d8f1d3e,
32'hbcc7035e,
32'hbcb1322c,
32'hbd0369bf,
32'hbcfe3715,
32'h3de4eec9,
32'h3ce71e8f,
32'hbb682596,
32'hbd56355b,
32'h3ce7186f,
32'hbc73ec8d,
32'h3d219f18,
32'h3b90d5c9,
32'hbc4465f3,
32'h3d201d52,
32'h3d7ced07,
32'hbc5f1592,
32'hbd34666c,
32'h3d31ceb8,
32'h3d3bb19a,
32'hbdb0f264,
32'hbd203717,
32'hbcc8c3d1,
32'h3d6912d7,
32'h3d2b07d2,
32'hbd791259,
32'h3cc423ff,
32'hbd8cde58,
32'hbcbfd288,
32'h3d90a917,
32'h3d3b399a,
32'h3db12b8f,
32'h3d1a1867,
32'hbc0f6e0f,
32'h3d2e2863,
32'h3c42aaa1,
32'h3c8942dd,
32'h3c48c3f3,
32'hbd994b2b,
32'h3cb1b957,
32'hbd3e0e6f,
32'h3ca6239a,
32'h3b78ea6f,
32'hbd6e6a1e,
32'hbd076574,
32'hbd439329,
32'hbc46d282,
32'h3cbf05da,
32'h3c230ce3,
32'h3da3f4c0,
32'h3d63784c,
32'h3dcbf438,
32'hbc751ca4,
32'hbbed3333,
32'h3db8b5f8,
32'hbd0c1dfe,
32'hbd3cc708,
32'h3ca5343e,
32'hbd9dc4ba,
32'hbd13c7c3,
32'h3f2a8c57,
32'hbf449159,
32'h3cdebe61,
32'h3ee8970b,
32'hbeabd3e7,
32'hbf1cfef5,
32'hbf2402a6,
32'h38ac719f,
32'hbddc80d0,
32'h3d08fdc1,
32'hbd7920ca,
32'hbda1d73b,
32'hbd8fe423,
32'h3e5ed5ef,
32'h3f082ee5,
32'hbe403d88,
32'hbeb96455,
32'h3e0b3f2e,
32'h3e238fdc,
32'h3dc91a7e,
32'hbf190442,
32'h3d0fdc9d,
32'h3f2c3447,
32'hbed52706,
32'hbef404e2,
32'hbe8704dd,
32'h3d2f03f7,
32'hbdbafc97,
32'h3e97b39e,
32'hbe32153a,
32'hbea1eeaf,
32'hbf0f6e03,
32'hbea251fc,
32'h3edc8c07,
32'hbf31ca56,
32'hbf04e74e,
32'h3e938db2,
32'h3c9556e0,
32'h3c19d987,
32'h3cd441fb,
32'hbdb68f2d,
32'hbec0894d,
32'hbdf4a5b3,
32'h3eedb915,
32'h3db1576d,
32'hbebc2001,
32'hbf07ef1d,
32'hbf4e0f00,
32'h3df94e51,
32'hbefe057d,
32'hbf003d98,
32'hbd350c0e,
32'h3f6c1c59,
32'h3d672026,
32'hbfab3c1f,
32'hbf03342b,
32'hbe6798e3,
32'hbe2e4f8e,
32'h3e583eff,
32'hbeccbcc2,
32'hbe608bd7,
32'hbec99621,
32'hbea6f35a,
32'h3ecbff63,
32'hbe24d063,
32'hbeac9c4d,
32'h3f3b292d,
32'hbecddb07,
32'h3e432172,
32'hbd006c06,
32'hbd020ff9,
32'hbf1c1b01,
32'hbc837799,
32'h3ea8c24f,
32'hbe646a0b,
32'hbe022d4f,
32'h3d48cf45,
32'hbedd448b,
32'h3e5724e8,
32'hbf0c1865,
32'hbe88c2d5,
32'h3d671f5b,
32'h3e5250f3,
32'hbd8dfd36,
32'hbf3ce0c2,
32'hbed05288,
32'hbeb56895,
32'hbd85fe2d,
32'h3e053c65,
32'hbf57a588,
32'h3e235ca9,
32'hbd320539,
32'hbe52de85,
32'h3f3ea8e5,
32'h3f3b2354,
32'hbf81667d,
32'h3f6d0adf,
32'h3ea3a43e,
32'h3e5824c0,
32'h3c6bec75,
32'h3c3220a4,
32'hbff294be,
32'h3d943277,
32'h3eb0e042,
32'hbdecf87c,
32'hbec729a0,
32'h3e5c7b36,
32'h3eb15697,
32'hbc4ba3a2,
32'hbfac418b,
32'h3ec70b71,
32'h3c26c1f2,
32'hbe9a8a28,
32'h3c7c1eb4,
32'h3f3e5f18,
32'h3eae4bf3,
32'hbe66e486,
32'h3d38ec1f,
32'hbec55c9c,
32'hbf8014f2,
32'h3ea25666,
32'h3e0cd121,
32'hbefabdc4,
32'hbd969ccf,
32'hbebe2810,
32'h3c91cb7b,
32'h3ed591d9,
32'h3e505add,
32'h3e9bfc8a,
32'hbd086d24,
32'hbda573a6,
32'hbfa5bedb,
32'hbe3b7634,
32'h3f479272,
32'h3e280289,
32'hbf830505,
32'h3f6f31fb,
32'h3ed2b6f4,
32'hbef9a8a4,
32'hbf3e8376,
32'h3ea9f3b9,
32'h3c4c8ba0,
32'h3e363a7e,
32'h3ee4785e,
32'h3f335e84,
32'h3e831944,
32'hbf5a7c7c,
32'hbe87b1ae,
32'hbf6ece4e,
32'hbed4aadf,
32'h3ecdab49,
32'h3ea8b368,
32'hbfa7ccea,
32'hbeaaf1fc,
32'hbf01df5c,
32'h3e24799f,
32'hbe95ac75,
32'hbf6be9ff,
32'hbdfd2b33,
32'h3d388cb1,
32'h3ca2abe2,
32'hbf11bcc9,
32'hbf0aa7f0,
32'h3ee3653e,
32'h3e84c5a5,
32'hbf3be395,
32'h3d04858b,
32'h3fa8fdd2,
32'hbf8da8bb,
32'hbf78cbc6,
32'h3f01c8cb,
32'h3dc50c27,
32'h3f096b53,
32'hbe7b6871,
32'hbe18e95f,
32'h3e1491a8,
32'hbe91f2a0,
32'hbeed87e3,
32'hbfdcad34,
32'hbe867152,
32'h3c103f1b,
32'h3f15033d,
32'hbfa1d73c,
32'h3f26f0a6,
32'h3f01d2a4,
32'hbd70460a,
32'hbe4aebf4,
32'hbf4bb764,
32'h3d72f674,
32'h3c20f1ca,
32'h3d80a904,
32'hbf06fa51,
32'hbebaa648,
32'h3eb68d00,
32'h3e11d987,
32'hbe3e9345,
32'hbe94c5f7,
32'h3ef80665,
32'hbe91eddd,
32'hbf3af38f,
32'h3f1e5e39,
32'h3e9e9c6f,
32'h3ece046b,
32'h3eacd935,
32'hbf55f830,
32'h3e13c36f,
32'hbeb6da8a,
32'hbd8f0067,
32'hbfc58e42,
32'hbea34ba9,
32'h3db6e257,
32'h3c34924f,
32'hbefa0317,
32'h3f84909f,
32'h3edf17d0,
32'hbe49198c,
32'h3f107bfa,
32'h3e326548,
32'hbf010bbf,
32'h3bf3f6ca,
32'hbda2727f,
32'hbf0d2bd2,
32'hbf0a6976,
32'hbf3afc7c,
32'hbdb71f09,
32'hbf3a9e2b,
32'hbf818e51,
32'h3b9cb189,
32'hbe11ea07,
32'hbf0a4c59,
32'h3f0b3db7,
32'h3e10367e,
32'h3f1baf55,
32'h3ee03f92,
32'hbf4af6d6,
32'h3f25f654,
32'hbe98eb46,
32'hbe97ef3a,
32'hbf689dee,
32'hbf576294,
32'hbe09d033,
32'hbe8dd3e1,
32'hbf0d8254,
32'h3e50b7c1,
32'hbf24ad97,
32'h3e30df2d,
32'h3f40595d,
32'h3e2b8f5f,
32'hbfa5ac49,
32'hbd83e018,
32'hbd96510b,
32'hbefebe68,
32'hbe75097e,
32'hbea178af,
32'hbe4904f5,
32'hbf32f752,
32'hbee2ee7c,
32'h3ea49569,
32'h3d76e9b5,
32'hbf66cc68,
32'h3f24d50f,
32'h3e18fa81,
32'h3ef7ee07,
32'hbe07c9c4,
32'hbf19464e,
32'h3ec67cf2,
32'h3d40a9a4,
32'hbdbfd10a,
32'hc01bda1e,
32'h3f38f977,
32'h3eb82bd1,
32'h3f5cbb6a,
32'hbfb74021,
32'h3ef90eb8,
32'h3ee863a7,
32'h3f08e2e5,
32'h3f146856,
32'hbdaa0a60,
32'hbf343495,
32'hbd1bd376,
32'h39bb40eb,
32'hbfa9a76a,
32'hbdebc7b1,
32'hbeac471a,
32'hbe66c06c,
32'hbde9ab65,
32'hbf04b704,
32'h3ecb5e53,
32'hbe26d91e,
32'hbf6da993,
32'h3f143976,
32'h3dcf59a8,
32'h3f14c286,
32'hbd83e8b6,
32'h3eb0693d,
32'h3f1f14af,
32'h3f2818f9,
32'h3f120b68,
32'hbf169c4f,
32'hbc8b4360,
32'h3e844f51,
32'h3f1d1f5a,
32'hbf815a77,
32'h3eb2b060,
32'hbec6f8cd,
32'hbf713156,
32'h3daaf336,
32'hbefd3a32,
32'hbf9da424,
32'hbd7ff47a,
32'h3d4838e6,
32'hbf98b9e8,
32'hbecb61b4,
32'h3e9cffd1,
32'h3ed563e5,
32'hbecbb412,
32'hbf284525,
32'h3f10c2c6,
32'hbf593c7f,
32'hbf7bd689,
32'h3e8fc032,
32'hbda23ce2,
32'h3ef70c81,
32'h3edf91b2,
32'h3c784eb1,
32'h3e90b34c,
32'hbebb5df2,
32'h3e38b7c2,
32'hbf25d5e1,
32'hbeea2540,
32'h3e9d483a,
32'h3e9389c5,
32'hbf837d02,
32'h3ec7b6a9,
32'hbdb7dbed,
32'hbf9af459,
32'hbd57cc27,
32'hbf9f6e47,
32'hbf338108,
32'h3b54f7f5,
32'hbd8719bd,
32'hbe714a77,
32'hbef0ec94,
32'hbe41c542,
32'h3c3f3f60,
32'hbda75398,
32'hbfab0c5d,
32'h3d7f27c2,
32'hbed8085b,
32'hbf8d5258,
32'h3ee4c66c,
32'h3e7a9e4f,
32'h3f7d479a,
32'hbd5ce8f2,
32'hbe9294b4,
32'h3f058732,
32'hbeeea4af,
32'h3eb99c05,
32'h3c0116ce,
32'h3f14238f,
32'h3e72d198,
32'h3dfbae29,
32'hbf5bed43,
32'h3e664ccf,
32'hbee51573,
32'hbf3694ff,
32'h3e9a1fc0,
32'h3e81e454,
32'h3e31c8fc,
32'hbd1a075e,
32'h3c687a65,
32'hbf4dc122,
32'hbe414da5,
32'hbf7c1b90,
32'hbe20cd24,
32'hbea64b91,
32'hbf41c6d5,
32'h3e954203,
32'hbe88da55,
32'hbf8f2fc3,
32'hbcb3d710,
32'h3e2611ed,
32'h3e8922b9,
32'h3e16c67b,
32'h3e8ea388,
32'hbdcf16a4,
32'h3f028acc,
32'h3f0973f3,
32'hbf53f0c2,
32'h3edcbae8,
32'h3bf3af64,
32'hbf004096,
32'hbfcaf12e,
32'hbec8b237,
32'hbf6fa082,
32'h3f070957,
32'h3dad1d5f,
32'hbed5b03a,
32'hbee51fc2,
32'hbda33a61,
32'h3ceb5f51,
32'hbf0eec78,
32'hbd85ca00,
32'hbf81dbb9,
32'h3e724f1f,
32'hbedd3186,
32'hbf6781b8,
32'h3e40cc47,
32'hbe7ac610,
32'hbfa10a90,
32'hbe03ce01,
32'h3dadbab4,
32'h3efe36ac,
32'hbe7e5fed,
32'h3de991cc,
32'hbe612230,
32'h3ebe869e,
32'h3f07be0f,
32'hbf4dc555,
32'h3ebc1af1,
32'hbe6fee19,
32'h3ddf1f97,
32'hbfb4bab1,
32'h3d181da2,
32'hbf1f72d1,
32'h3f2eb411,
32'h3e198679,
32'hbe8cf13c,
32'hbe13b4a4,
32'hbd801da7,
32'hbd6ebfa3,
32'hbf31d5f1,
32'hbe1c626c,
32'hbf810a10,
32'hbe3a1b2e,
32'hbed8f982,
32'hbfa87638,
32'h3e1fffee,
32'hbf8bfc6d,
32'hbf348b52,
32'hbd2bdf47,
32'h3d272e4a,
32'h3f0d2cae,
32'h3e4b9e2c,
32'h3f828b14,
32'h3e75f64a,
32'h3e600f3d,
32'h3e50033b,
32'hbfc129e8,
32'h3ea2da78,
32'h3fbdce1d,
32'h3f30c7e2,
32'h3ea4c46c,
32'hbf9a67d9,
32'h3eccd457,
32'h3f0ebbfc,
32'h3d64821c,
32'hbe82e867,
32'hbe55dcbc,
32'hbd3d6129,
32'h3bd73a66,
32'hbe6e4d50,
32'hbe4ffea4,
32'hbd3f2a4d,
32'hbf21ec6a,
32'h3d365e56,
32'hbf2c1e65,
32'hbd948636,
32'hbf7478bb,
32'hbf8a8027,
32'hbe868ae7,
32'h3de71960,
32'h3e2fb452,
32'h3cf78f4e,
32'h3f6ada2e,
32'h3e9fa16d,
32'h3e9de5b1,
32'hbeb5a690,
32'hc00841f3,
32'hbc5b9e80,
32'hbf07e872,
32'hbde60620,
32'hbf716c9e,
32'h3ea432b2,
32'h3e0ed794,
32'h3f82bfc6,
32'hbe54d9bd,
32'hbe60902c,
32'hbefc97af,
32'hbd708464,
32'hbcdba1ca,
32'hbe3b366e,
32'hbe209f8c,
32'hbf031504,
32'h3eb8f3ba,
32'hbdfa3a08,
32'hbf603368,
32'h3e2c679f,
32'hbe03c224,
32'hbf9ecdd6,
32'hbe32652a,
32'h3b045cf4,
32'hbe9503fe,
32'hbf029976,
32'hbe61139f,
32'h3ec31dd3,
32'hbeb9c16e,
32'hbf16df78,
32'hc0076dea,
32'hbce051b3,
32'hbe819c50,
32'hbf893658,
32'hbf24c4b0,
32'h3f5c1b09,
32'h3d11db8a,
32'h3f2532a0,
32'h3f5d4f0b,
32'hbf2ea616,
32'hbd24323a,
32'hbd513dcc,
32'hbdc365b9,
32'hbf2e602a,
32'hbdafa623,
32'hbe48ddf5,
32'h3e887d24,
32'hbdbf287b,
32'hbfb95531,
32'h3f196ff1,
32'hbf2e4b92,
32'hbfd81ac7,
32'h3e9fbcc0,
32'h3bebaef4,
32'hbf201b4d,
32'hbf318a53,
32'h3dc3ac5f,
32'h3e457607,
32'h3f431a61,
32'hbda22b33,
32'hbfb1f7bb,
32'h3cab05f4,
32'h3e829a17,
32'hbec2f976,
32'h3d93db11,
32'h3ef097e8,
32'hbd723395,
32'h3f5027f8,
32'h3f597138,
32'hbe5a977d,
32'h3cf1a10a,
32'hbcb1c1e8,
32'hbc132da6,
32'h3e7b4b67,
32'hbea59dcf,
32'hbe479adb,
32'hbf00639b,
32'hbd90fa04,
32'hbf879aec,
32'hbd284d76,
32'hbf903abc,
32'hbfd0c0b5,
32'h3f23fe80,
32'hbcd4e701,
32'hbcb2b056,
32'hbdf1a88f,
32'h3ef9bbca,
32'h3f128600,
32'h3ea3582b,
32'hbca2c398,
32'hbf6ff93a,
32'hbdaa8d6a,
32'h3f892f2a,
32'h3c9ad73a,
32'h3e189065,
32'hbf4e016b,
32'hbdedd8a7,
32'h3b92a8ff,
32'h3f2503eb,
32'h3acd3946,
32'hbda3350d,
32'h3d81ada0,
32'h3d3847e8,
32'h3e7f2f35,
32'h3c7ee010,
32'h3de2b552,
32'h3b9fc15e,
32'hbbd8fd5b,
32'hbf3bd2b2,
32'h3efc9eaf,
32'hbe23ce8c,
32'hbf823c53,
32'hbdc5a393,
32'hbd40178c,
32'hbe561e07,
32'hbda36c26,
32'h3ebe1907,
32'h3f0f7df5,
32'h3f0f746f,
32'hbd583c9c,
32'hbf248862,
32'h3c777cd8,
32'hbe78ec17,
32'hbc74de7e,
32'hbbaae9bd,
32'h3e868cae,
32'h3b81682c,
32'hbcc8a5e6,
32'hbdb01e80,
32'h3de9c6e6,
32'hbd04d180,
32'hbd38127f,
32'hbdbe0601,
32'h3ea8d967,
32'h3d5f4dbb,
32'hbd261f0a,
32'h3f2a36b8,
32'h3c0937d8,
32'hbd42fb64,
32'h3f233233,
32'h3e92f0b8,
32'h3e242f66,
32'hbeef3ded,
32'hbce1551c,
32'hbf1ed5ee,
32'h3dd171f7,
32'hbec4a37d,
32'hbca9db51,
32'h3d1b6ae9,
32'h3b829554,
32'hbe0bf3c8,
32'hbdb821d0,
32'hbda73bb3,
32'h3d8a4e8d,
32'hbd8af4d3,
32'h3bf07204,
32'hbe2ddadd,
32'hbdaf3813,
32'hbd4570bf,
32'hbcbe6206,
32'h3c84e289,
32'h3b07facd,
32'hbcad7034,
32'h3d01183e,
32'hbd236214,
32'hbd03e00e,
32'h3ca6b3d2,
32'h3bdb632e,
32'hbdb44562,
32'h3d90ebfa,
32'hbd7cd23e,
32'h3b6b5499,
32'h3d87e193,
32'h3da1d896,
32'hbc84658c,
32'hbd6c4914,
32'h3c4a2e7f,
32'hbb976a68,
32'h3dd4fd0a,
32'h3c1e8a38,
32'hbc307563,
32'h3c3f708f,
32'h3ce99a2a,
32'h3c37799b,
32'hbdeb0ac8,
32'h3d0f1940,
32'hbd09a36c,
32'h3d578126,
32'h3cc00074,
32'hbb2ab8dd,
32'h3cb9b2a5,
32'hba4245f9,
32'h3d76db8d,
32'hbda8a077,
32'hbca3e40c,
32'h3d049553,
32'h3ce19e16,
32'hbd1c6b84,
32'hbd1c6239,
32'h3cb59af5,
32'h3d0a9cfc,
32'hbc2fced6,
32'hbd8d70c0,
32'hbdd86013,
32'h3d77b9a8,
32'hbd362569,
32'hbd1eaccc,
32'hbd8e6d66,
32'hbccaea58,
32'hbd678ead,
32'hbb2f3ba3,
32'h3b244cea,
32'h3bb0277c,
32'h3d3c3ad4,
32'h3c09341d,
32'hbcd308f8,
32'hbd32090d,
32'hb978a3a4,
32'hbc2f8edd,
32'h3d3178d3,
32'h3ce9669a,
32'h3d1ffe55,
32'hbc87a4ba,
32'h3d93d986,
32'h3d38adca,
32'h3ca09bdb,
32'hbb90924f,
32'h3caf74e8,
32'hbd38ead2,
32'h3d95da74,
32'hbcbbd143,
32'h3c7c3940,
32'hbc5d728d,
32'hbd3d0775,
32'h3d01d96f,
32'hbd66230f,
32'h3c8e0581,
32'hbcc11ea3,
32'h3d106d63,
32'hbd8105dc,
32'hbd65c006,
32'hbd9753d6,
32'h3d846f6e,
32'hbd46fde7,
32'h3dbfda3f,
32'h3d287619,
32'h3dcc636b,
32'hbcd64c69,
32'h3b935c7b,
32'hbda42d29,
32'hbce2a213,
32'hbd1f9023,
32'h3d2092de,
32'hbdc33104,
32'hbd40efdb,
32'hbd57e8c5,
32'hbca8369f,
32'h3d261e68,
32'h3d49f911,
32'h3b5e5843,
32'h3cffbe15,
32'hbd3757d6,
32'h3d36a540,
32'hbcf8831d,
32'h3db4d650,
32'hbd849acc,
32'hbda96895,
32'hbc12b14a,
32'h3d5bda24,
32'hbbec78c4,
32'hbbd8660b,
32'h3d497297,
32'hbd393637,
32'hbc2b4f0f,
32'h3daadd4b,
32'hbcc95da3,
32'hbd7dfeb4,
32'h3c4083fd,
32'hbc526d59,
32'h3d814fa4,
32'hbda52275,
32'h3d055aaa,
32'h3d785664,
32'hbd167156,
32'h3d462431,
32'h3ce2aa48,
32'hbc0366fa,
32'h3d4d53f6,
32'hbde1465a,
32'h3c7f2eb1,
32'h3cc627ac,
32'h3dc2c6d0,
32'h3dda85cb,
32'h3ddcb456,
32'h3d3a7660,
32'h3d877be4,
32'h3be4fc10,
32'hbd1e064f,
32'h3db72938,
32'hbd78fad5,
32'h3da59c7f,
32'hbca2016d,
32'hbd865aed,
32'hbc59193b,
32'hbd39b8c5,
32'hbccf87fd,
32'hbde090d0,
32'h3db1ca6c,
32'h3ca7a364,
32'h3d57b043,
32'h3cd54be9,
32'h3dcee566,
32'hbd48d3c6,
32'h3d2af223,
32'hbdabf5a2,
32'h3ccc2992,
32'hbc9fcb22,
32'hbd84ac84,
32'hbd545a2d,
32'h3da2b556,
32'hbbc7bbf3,
32'h3c62375c,
32'h3c9f3f05,
32'hbd075eaa,
32'hbc300200,
32'h3d199500,
32'hbda2bd7d,
32'hbca60176,
32'hbd22f6a3,
32'hbb195d9d,
32'h3c6dc94f,
32'hbcfbcef9,
32'hbddc1c56,
32'h3deae9cd,
32'hbd50cf06,
32'hbdbc3d53,
32'hbcee1369,
32'h3cddf874,
32'h3d1946eb,
32'h3d8bf272,
32'hbcad558b,
32'hbd22c2f5,
32'h3c678dc0,
32'h3c0be11e,
32'h3d975ec6,
32'h3c8dac8f,
32'hbd9231b3,
32'hbce63a94,
32'h3d2fdb34,
32'h3dae5246,
32'hbd07261d,
32'hbbc4b7b3,
32'h3d2742b0,
32'h3d3cd551,
32'h3c73ac90,
32'h3cd6a33e,
32'hbdcf6d20,
32'hbc998bb6,
32'hbce02e84,
32'hbd2f61e8,
32'hb92403b4,
32'hbd90bb40,
32'h3d5371cd,
32'h3e06e0b8,
32'h3d599202,
32'h3edd1948,
32'hbe140f83,
32'h3d3f9853,
32'h3d62ce2b,
32'h3dd4e983,
32'h3c806a42,
32'hbd2fd4f9,
32'h3d09e813,
32'h3d9ed9cb,
32'h3d83fda4,
32'h3e44fdb0,
32'hbe987fd8,
32'h3bc2316c,
32'hbcd6b307,
32'h3e15a2ef,
32'h3d13a1f3,
32'hbc826cf0,
32'hbe52dec4,
32'h3d5107e3,
32'hbf3dff6e,
32'hbb94857c,
32'h3f4cb11b,
32'hbe2e9508,
32'h3e9ff273,
32'h3c99b08a,
32'hbd784650,
32'hbe2d741b,
32'h3f54cb34,
32'h3e221296,
32'hbb31a7e9,
32'h3f4eef70,
32'hbd59488e,
32'hbddab86b,
32'hbdc6e6fc,
32'h3daab1dd,
32'h3e3f2dda,
32'h3db55d31,
32'hbd98f450,
32'hbd1c0e7a,
32'hbd2cfff5,
32'h3e929a8b,
32'hbf20127e,
32'h3cf08d2f,
32'hbc5abcfd,
32'h3f37b768,
32'h3ee77c1a,
32'hbe23657f,
32'hbefcc183,
32'hbda1dd65,
32'hbf4739a7,
32'h3c284f87,
32'h3f734b71,
32'hbebf50e5,
32'h3e937d89,
32'hbd9de9bf,
32'hbe2a3218,
32'hbbec95a4,
32'h3f1b0abf,
32'h3dbd4614,
32'hbe7f3645,
32'h3ec2b75b,
32'hbe00e927,
32'hbe854a87,
32'h3ca71841,
32'h3d11a2b3,
32'h3e0cb222,
32'hbda68fa5,
32'h3dc83b75,
32'hbc4d41bf,
32'hbd99cd53,
32'h3e897e00,
32'hbebf935b,
32'hbd33c336,
32'hbec05765,
32'h3e209c11,
32'h3ddad7e2,
32'hbfac1326,
32'h3dd12ea2,
32'h3c4f7eb4,
32'hbe8cfebe,
32'hbdb3dc0c,
32'h3f0b3fb6,
32'h3d179dea,
32'h3def83f4,
32'h3c1e5843,
32'hbf1cbb23,
32'hbcb89075,
32'h3f1b4912,
32'h3e379ff8,
32'hbe11b1da,
32'h3e4c018c,
32'hbd8b7de3,
32'hbee3de16,
32'hbc2622f6,
32'hbd5fbbfd,
32'h3de06a7d,
32'hbcbf6d84,
32'h3cc55a96,
32'hbd8d1b4f,
32'hbd5eca1e,
32'h3e459e2e,
32'hbe80368b,
32'h3d431965,
32'hbed73d90,
32'hbe0a1282,
32'hbe20b1bc,
32'hbfb440c0,
32'h3e469a4f,
32'h3d69197b,
32'h3ead0f9e,
32'hbd0c2172,
32'h3e409ed8,
32'h3e3f01d4,
32'h3e641018,
32'h3d99c843,
32'hbf392107,
32'hbc555ac8,
32'h3f2e99b2,
32'h3e628299,
32'hbc11b57e,
32'hbe1962b0,
32'h3dbaf50a,
32'hbed2b617,
32'h3d7f877c,
32'hbc8f1dd4,
32'h3ea3cf62,
32'h3ce92dff,
32'h3c87d61d,
32'h3d264bc9,
32'h3d1654e2,
32'hbd8cd8c8,
32'hbec15084,
32'hbd18483d,
32'hbee72708,
32'h3d36fd16,
32'h3e3a307d,
32'hbfb6b2f9,
32'h3de5e768,
32'hbd90b4f3,
32'h3eba2f31,
32'hbca5d5a2,
32'h3e0f5151,
32'h3e6181e4,
32'h3e3921ea,
32'hbc66128d,
32'hbf5994b3,
32'h3f09295e,
32'h3f784eb2,
32'h3f26a6c4,
32'hbe116fab,
32'hbd99b612,
32'hbcc4106b,
32'h3d19393f,
32'h3eed1edf,
32'hbe2ee88c,
32'h3eacd4d9,
32'h3c5b0195,
32'h3dd03f15,
32'h3dae748f,
32'hbdc85832,
32'hbe6a8c3c,
32'h3e5217dd,
32'hbab6819b,
32'hbee79589,
32'h3e6345ff,
32'h3e8dac84,
32'hbfa69656,
32'hbf4a2899,
32'hbbb515fe,
32'hbd9d33a9,
32'hbdd3f0a7,
32'h3e335576,
32'hbe669e46,
32'hbe365b25,
32'h3a44baeb,
32'hbf5e37eb,
32'h3e090c33,
32'h3e169a8e,
32'h3f433eda,
32'hbdd509ed,
32'h3f0980ab,
32'h3e83aae1,
32'hbe0fdc22,
32'h3f1713ae,
32'h3d66ef51,
32'h3e85a270,
32'hbc601334,
32'hbd18cc97,
32'h3dfc3bc2,
32'hbd3161d9,
32'hbe8ecbd1,
32'h3e408638,
32'h3c74fadb,
32'hbe76ed68,
32'h3ec3f7e5,
32'h3d8be393,
32'hbf61730f,
32'h3e42a36f,
32'h3d838cf1,
32'hbf4acb3b,
32'hbe784c2a,
32'h3f4b7465,
32'hbdf37c72,
32'hbe70a239,
32'hba825e3d,
32'hbf11d661,
32'h3e07f9ec,
32'hbe8f2f9b,
32'h3f5a06b4,
32'hbe044bb3,
32'h3f430af3,
32'h3e0a45be,
32'hbecb6ac8,
32'hbed2a024,
32'hbf24d445,
32'h3e9b3aec,
32'hbdac5703,
32'h3c308c14,
32'h3db28274,
32'hbdf289ef,
32'hbee527bf,
32'h3e83c181,
32'hbd132ff2,
32'hbed139cd,
32'h3c9defe9,
32'hbe06564c,
32'hbf7cf2ba,
32'h3e777b85,
32'h3da4feb0,
32'h3e93365e,
32'hbea95ba7,
32'h3cbfe483,
32'h3cc9e552,
32'hbe816c8c,
32'hbdc1cf29,
32'hbee45a18,
32'h3df19e52,
32'h3f12f9b8,
32'h3ee16bf6,
32'h3c40c213,
32'h3e318f37,
32'h3e867cd4,
32'hbe81d6aa,
32'hbd56d3d5,
32'hbf133263,
32'h3eca9a94,
32'hbd6f2ecf,
32'hbcd04e83,
32'h3e394d77,
32'hbd88b8e3,
32'hbe732b5b,
32'hbeb79b29,
32'h3cc323c8,
32'hbec6d80e,
32'h3e924fb5,
32'h3f132358,
32'hbf5166b5,
32'h3e017420,
32'h3cdb5776,
32'h3b912007,
32'hbea92b49,
32'h3ef8340e,
32'hbe1db276,
32'hbdd0fd92,
32'h3cc857e7,
32'hbf41dd96,
32'h3e9d6315,
32'h3ec8a25e,
32'h3eaecdc3,
32'hbe1aacae,
32'h3ed8e809,
32'h3e653c6e,
32'hbde1bdab,
32'h3e642cd8,
32'hbf2865c1,
32'h3e539f58,
32'h3bd0e42c,
32'h3b92d360,
32'hbd5a6109,
32'hbb5458d6,
32'h3ce0a2ab,
32'hbeb6e030,
32'hbe988844,
32'hbeeca5d0,
32'h3f285c40,
32'h3f813e36,
32'hbfb6326d,
32'h3ec764cc,
32'hbd83637c,
32'hbdef0dfb,
32'hbee88694,
32'h3eaac66e,
32'hbcee70d4,
32'h3d356567,
32'hbc51d66e,
32'hbf71568d,
32'h3f2775a6,
32'h3ed0ea78,
32'h3e4fa22b,
32'hbea2d649,
32'hbd885711,
32'h3e1caf55,
32'hbee61adf,
32'hbed66352,
32'hbef8df28,
32'h3e85e6e0,
32'hbd32a3e0,
32'h3baecbea,
32'hbe2e1da4,
32'hbc98b3a7,
32'hbea24ea7,
32'hbd10f134,
32'hbe1be99f,
32'hbf04065c,
32'h3f39b5df,
32'h3f86be7f,
32'hc00c34cc,
32'h3f459374,
32'h3d81882a,
32'hbe0bb924,
32'hbeae150c,
32'hbeb01506,
32'h3ecd49ea,
32'h3e04c8de,
32'h3c826d86,
32'hbfd9cb6d,
32'h3ddd0e14,
32'hbe932e92,
32'h3d40e927,
32'hbe71faf4,
32'hbe6749b0,
32'h3f3b63ea,
32'hbe62030b,
32'hbf5268d1,
32'hbee25b37,
32'h3e173fe4,
32'h3c851b1c,
32'h3da6d1d1,
32'hbe0c358e,
32'h3ce7da76,
32'hbdac3e92,
32'h3f529ac1,
32'hbd5e4af0,
32'hbd385620,
32'h3f2c086c,
32'hbef3b734,
32'hbe28b9bf,
32'h3ee68af6,
32'h3d8648fe,
32'hbd567851,
32'hbe8a6089,
32'hbf2dae08,
32'h3f61b8fb,
32'hbe1f3664,
32'hbd63e2da,
32'hbf220e45,
32'h3bfc18dd,
32'h3ed3e5b7,
32'h3e0d1249,
32'hbe5fff76,
32'h3dae5b10,
32'hbe4bb84e,
32'h3d7c9bab,
32'h3e144c82,
32'hbe28bdb9,
32'h3e99c994,
32'hbc8a0e77,
32'hbd93cfe6,
32'hbdd1fea6,
32'h3d00927b,
32'h3e41f84e,
32'h3f1e5125,
32'hbc34f3d1,
32'hbf10c930,
32'h3e79cdb6,
32'h3f227136,
32'hbf05d4c1,
32'hbd96e9fc,
32'hbda42e34,
32'hbdb5255d,
32'h3e1d92d8,
32'h3f500003,
32'hbeea9622,
32'hbdaf2446,
32'h3b454465,
32'hbdd5b67a,
32'h3e3a6677,
32'h3ef5fa3c,
32'hbe1d4137,
32'h3e955cb9,
32'hbe48ed4d,
32'h3dfcd7ae,
32'hbe7f8c3d,
32'hbe3de8c8,
32'hbeea5889,
32'h3ea6fda2,
32'hbcb8b7bc,
32'h3cced1df,
32'hbe0b2a50,
32'h3b850006,
32'h3f057948,
32'h3e4070cf,
32'hbe13e065,
32'hbf0478cf,
32'h3f83c35c,
32'h3e9e05dc,
32'hbe3cdd85,
32'hbebc38b8,
32'h3d4ce0ef,
32'hbea983c9,
32'hbe5dbb76,
32'h3ea6a89a,
32'hbe515b6a,
32'hbef50cae,
32'h3ddba052,
32'hbf6e109f,
32'h3e88e5e3,
32'h3f7dd934,
32'h3d11c662,
32'h3eb52654,
32'hbe6d57de,
32'hbca6d9b8,
32'hbeadf757,
32'hbe67855f,
32'hbe796dc9,
32'hbe4a7c93,
32'hbdb8c625,
32'hbd13a857,
32'hbe4bcb45,
32'hbca069ed,
32'hbe296dce,
32'hbe41a557,
32'h3c83b8b7,
32'hbe93da0b,
32'h3f8f748d,
32'hbdf8156c,
32'hbe8552ee,
32'h3cb05977,
32'h3d0ed78f,
32'h3e974569,
32'h3e34d3d0,
32'h3d085150,
32'hbea8182e,
32'hbf383b29,
32'h3d59cfaa,
32'hbf6c191e,
32'h3e64b2e9,
32'h3f00431b,
32'h3cf28123,
32'h3eacb22e,
32'hbe58b60c,
32'h3cc4d05a,
32'hbbedf747,
32'hbd24f220,
32'hbdf711fe,
32'h3e0ca496,
32'hbc12f3c8,
32'h3c3181b3,
32'hbe07364f,
32'hbb0611bf,
32'h3bdcbefa,
32'hbe45a9b0,
32'hbde68564,
32'hbecdc65a,
32'h3db5842f,
32'hbe40bf63,
32'hbf43022f,
32'hbdeaa87f,
32'h3d739aad,
32'h3ed893af,
32'hbf3bc62b,
32'hbcc1903f,
32'h3ea87531,
32'h3ecabdd2,
32'h3caf1bff,
32'hbedc7355,
32'hbd22e516,
32'h3e219a9e,
32'h3d03158a,
32'h3e57cf55,
32'hbd72874d,
32'h3d07b066,
32'h3dfe705f,
32'hbd914cc2,
32'hbe1ede34,
32'hbdd3215d,
32'h3c29fd80,
32'h3cbc0f76,
32'hbdf05ed6,
32'h3ce45a8a,
32'hbe503c67,
32'hbcbdbf68,
32'hbd1e9da3,
32'hbebf26b7,
32'h3d0974a5,
32'hbe6604ad,
32'hbe147761,
32'hbeda7ac5,
32'h3d9b8595,
32'h3edce0ac,
32'hbf35345d,
32'hbe1bd65d,
32'hbef8435d,
32'hbda47183,
32'hbba177dd,
32'h3c1e3c4c,
32'hbd5b67b6,
32'h3f43bd6d,
32'hbe46cc27,
32'h3e32d53f,
32'h3eab8d4f,
32'h3d5d0b63,
32'h3d97cf95,
32'h3eecfb87,
32'hbe1298d1,
32'hbc734171,
32'h3db6bdc0,
32'h3d0dc21a,
32'hbf3c28fa,
32'hbc343c97,
32'hbd4b6ec3,
32'hbed621cc,
32'h3de8faed,
32'hbf08add1,
32'h3eab2698,
32'hbd885644,
32'hbf806490,
32'hbf332a2b,
32'h3d461fa0,
32'hbdd06507,
32'hbec4c2ce,
32'hbe9785db,
32'hbf1c7d1b,
32'h3ef06361,
32'h3c102c73,
32'hbe8ddef2,
32'h3d5a4fe4,
32'h3edc3965,
32'hbe167f4a,
32'h3d5e4f3c,
32'hbcfb91f4,
32'hbd6fc103,
32'h3c866577,
32'hbd0624a4,
32'hbde73e5a,
32'hbc88cd4b,
32'h3cf7440c,
32'hbde5f13a,
32'hbdaaa2f7,
32'h3ca9b456,
32'h3d222465,
32'h3e3c1141,
32'hbd25f95e,
32'h3e9e0a9e,
32'h3e572450,
32'h3e100a0c,
32'hbc3708e9,
32'hbdd5bdfc,
32'hbc039650,
32'hbe77bc96,
32'hbeb96a12,
32'hbe93aa03,
32'hbdba39d8,
32'h3e2b5ccc,
32'hbca1c99b,
32'hbdbf2555,
32'h3c9630a6,
32'h3f069d09,
32'hbd46f654,
32'hbc608e68,
32'h3ea4e25b,
32'hbd7302f9,
32'h3d62c50c,
32'h3e4f01cd,
32'h3a1d2d10,
32'hbbe25fce,
32'hbdc39c14,
32'hbd81488c,
32'h3ccd4cb0,
32'hbd77b855,
32'hbcbe8cf4,
32'hbed215ab,
32'h3d659a87,
32'hbd72c444,
32'h3eb91bb7,
32'h3e0f83ea,
32'hbd97a563,
32'hbe0fed19,
32'h3be7d9e0,
32'hbef160f8,
32'h3d6c95c1,
32'h3ec9c6bb,
32'hbd9d8d41,
32'h3eee45e7,
32'hbc882877,
32'hbeca23db,
32'hbd78d7a8,
32'h3c641bf7,
32'h3cc57a12,
32'hbc68a478,
32'hbb949e74,
32'h3dd4232e,
32'h3d51ab3a,
32'hbc40bfe1,
32'h3cbeb8f1,
32'hbbf1885f,
32'h3c2b600a,
32'hbc0a3779,
32'hbd5795b1,
32'hbdc095e0,
32'h3d8bff70,
32'hbd80c4fd,
32'hbb77294e,
32'hbd105fb6,
32'hbcf3e922,
32'hbd598ba5,
32'h3d8a86af,
32'h3c596503,
32'hbce883ef,
32'h3d256832,
32'h3dc427d1,
32'h3dcc5257,
32'hbd2ff0aa,
32'h3babd8ef,
32'h3d26ab58,
32'h3b79cc07,
32'hbd2daa9a,
32'hbd56cbf2,
32'h3ddc0b43,
32'hbd397ac9,
32'h3c0601ae,
32'hbcfab8e6,
32'hbd868b68,
32'hbd8fe5cd,
32'h3bda40f5,
32'h3cf6a362,
32'h3d9235bf,
32'hbd1fea15,
32'h3d163005,
32'h3d1ec23a,
32'hbc5cb342,
32'h396145c3,
32'hbd00f8da,
32'hbd39b723,
32'h3d1fb638,
32'hbd2f09fb,
32'hbde46aa8,
32'hbbd107bc,
32'hbb841136,
32'hbce9296e,
32'h3de61bee,
32'hbd0b1369,
32'h3db3c021,
32'hbca0986d,
32'h3d7d50da,
32'hbd198006,
32'h3d93b674,
32'hbaefeac9,
32'hbc5fdcaa,
32'h3d31e46d,
32'hbd3c0f6a,
32'h3d0ccc60,
32'h3d9adfb6,
32'hbd312b6c,
32'hbd7120f4,
32'hbb42ae9b,
32'h3d3daea3,
32'h3dab0088,
32'hbd735aba,
32'h3d667f7c,
32'hbd659db5,
32'hbd642380,
32'h3c3900dc,
32'h3c9de3d3,
32'h3d945b31,
32'hbbb22bd9,
32'hbde830dd,
32'h3cb4498f,
32'hbd9381e0,
32'hbd37bb4f,
32'hbcab328f,
32'h3d6431c2,
32'h3d1e6e47,
32'h3bf23806,
32'hbd84c236,
32'h3d23543b,
32'hbd9c86e1,
32'h3d7c6faf,
32'h3b9f3baf,
32'hbd900ebb,
32'hba355598,
32'hbd43cb2f,
32'hbcd13634,
32'hbd0fc1e2,
32'h3dd9f273,
32'hbdad5bc1,
32'hbc3d1ee8,
32'hbd01d747,
32'h3d7c3992,
32'hbc66514a,
32'hbd5ce8d5,
32'h3cc76900,
32'h3d49fde7,
32'hbd57966a,
32'hbd202830,
32'hbd56ce81,
32'h3ca0a16a,
32'hbd4c40c4,
32'hbcf2ff73,
32'hbc6bcb48,
32'hbdd52812,
32'h3d462b10,
32'hbc802175,
32'h3ddaf18b,
32'hbd9445a5,
32'hbdad16d3
};
	assign weight = {ROM[addr],ROM[addr+1],ROM[addr+2],ROM[addr+3],ROM[addr+4],ROM[addr+5],
						ROM[addr+6],ROM[addr+7],ROM[addr+8],ROM[addr+9],ROM[addr+10],ROM[addr+11],
						ROM[addr+12],ROM[addr+13],ROM[addr+14],ROM[addr+15],ROM[addr+16],ROM[addr+17],
						ROM[addr+18],ROM[addr+19],ROM[addr+20],ROM[addr+21],ROM[addr+22],ROM[addr+23],
						ROM[addr+24],ROM[addr+25],ROM[addr+26],ROM[addr+27],ROM[addr+28],ROM[addr+29]};
endmodule 