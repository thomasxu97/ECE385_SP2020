module weight_mat_w1(
	input [14:0] addr,
	output [31:0] weight
);
	parameter ADDR_WIDTH = 15;
   parameter DATA_WIDTH = 32;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
32'hBCD6C54C,
32'h3D821705,
32'h3D317BF1,
32'hBCDD0DB5,
32'hBD88D9F1,
32'hBC463AF5,
32'hBD1E508C,
32'hBC22AC22,
32'hBD468956,
32'hBD7D7352,
32'hBC7F0974,
32'h3D631564,
32'h3D97A41A,
32'hBD4E33CC,
32'hBD833006,
32'h3CE94A1D,
32'hBD0180DE,
32'hBD3B8610,
32'hBD19378E,
32'h3C7C5FC3,
32'h3CA58C59,
32'hBD1F4833,
32'h3D03BF1F,
32'h2EDF5BA8,
32'h3C8CD1B0,
32'hBD9D7A36,
32'h3CE32247,
32'hBD85476B,
32'hBC137EA0,
32'hBC2C2F07,
32'h0ED61789,
32'h3CD1EC07,
32'hBC0F8FF9,
32'h3D53A11D,
32'h3D1590EC,
32'h3D541B33,
32'hBD9AEEC4,
32'hBD9A893A,
32'h175BC538,
32'hBD51BE02,
32'h1DF82973,
32'hBDB42158,
32'h3D9BFECE,
32'h3CFF9868,
32'h3DBA8035,
32'hBCA06F44,
32'h3DC20BB8,
32'h3CA1F580,
32'hBD6A5644,
32'h1DDC6646,
32'hBD9825F1,
32'hBCFD9974,
32'hBCA783A8,
32'hBD2D360D,
32'h3D84A97A,
32'hBCD2A216,
32'h3CBF45DA,
32'hBCE36A1D,
32'hBD1B94AC,
32'hBCD4B4CC,
32'h3DBECF72,
32'hBCCAFB28,
32'hBD30FAB0,
32'h3C85A312,
32'h3D75A0D3,
32'h3CFF1DF6,
32'hBD8F849B,
32'hBCA140CA,
32'h3C8C5EAE,
32'hBD97ABC4,
32'hBCE673A0,
32'h3D4AF724,
32'h3C85DBF3,
32'h3DB529F7,
32'h3D9A202F,
32'hBCE8F1E5,
32'h3D2C11C6,
32'hBC27F4BD,
32'hBC9A0244,
32'h3DE049EC,
32'hBC3CA6CF,
32'hBD98AC79,
32'h3D1A4AE1,
32'hBCE8C7E2,
32'h3C71E4F3,
32'h3D7417A1,
32'hBD583ADE,
32'h3D77F2A6,
32'h3CA7CE99,
32'h3D09C21C,
32'h3D65D628,
32'hBC9C954F,
32'h3D17F2B1,
32'h5DE2BCFB,
32'hBD396CDD,
32'h3D32FDDC,
32'hBDD07080,
32'h3DB99CB0,
32'h3C824154,
32'hBD90C993,
32'h3D33B079,
32'hBDBBF1F2,
32'hBC2E9691,
32'hBD7B5DCB,
32'hBD0DA511,
32'h3CCF553A,
32'hBD7C241B,
32'hBD837DAC,
32'h3DB9C065,
32'hBD1FBA45,
32'h3CA4D1CB,
32'hBC816F00,
32'hBC21CF4F,
32'h3D64BA0B,
32'h3D177D4F,
32'hBDAD3E96,
32'h3D1E3918,
32'h3D617B6D,
32'h3D7FDA77,
32'h3D608F16,
32'hBC9C714F,
32'h3D644A7E,
32'h3D7F2CD9,
32'h3CC35D65,
32'h3C99DA2A,
32'hBD19717C,
32'h3C8431AD,
32'h075CABEA,
32'hBD98D8DC,
32'hBC54207A,
32'hBCB5CF50,
32'hBDAC8193,
32'hBD9486E1,
32'hBD09F692,
32'hBC9D64DB,
32'h1DCC648E,
32'hBD412C64,
32'h3CBDE416,
32'h3D06E87B,
32'h3DBE1B49,
32'h1DCACF61,
32'h3C7B535D,
32'h3D2760B8,
32'h3D1211A8,
32'h5DF1511F,
32'hBDB989B2,
32'hBD27B3BB,
32'h3CF5F2EB,
32'hBD1B2545,
32'h3D5F9AF2,
32'hBD881115,
32'h3CBD435B,
32'hBCBE5691,
32'h3C0023CB,
32'h3D71AB47,
32'h3D6EF539,
32'h0EC82186,
32'hBD7530B0,
32'hBCCA41F1,
32'hBD92E122,
32'hBD8D0993,
32'hBD2F7DA9,
32'h3D8E1042,
32'hBD66732E,
32'h3D493954,
32'hBD3862DD,
32'hBD104C9A,
32'h3CC7FCAE,
32'h3C5CEF08,
32'h3C3D1225,
32'h3C80B1F5,
32'hBDCB99B4,
32'hBC895476,
32'hBD51A559,
32'h3CF8EF65,
32'h3C6E9847,
32'h3C5C3BC3,
32'h5DC5C4B2,
32'hBC65E19C,
32'hBD9AFF00,
32'hBD770B62,
32'h1DF935B9,
32'hBD429E58,
32'h5DC5DD1F,
32'h1DEDD544,
32'hBCC4E5EA,
32'h3D2F3C1B,
32'h2ED60A4F,
32'hBD98CC97,
32'h1DC1D593,
32'h1DCADA45,
32'hBD33A073,
32'hBD88AA27,
32'h17598C23,
32'h5DE9E670,
32'h3C8239BC,
32'h3CD2057B,
32'hBCB18EB4,
32'h2ECEC376,
32'h3DC6EFE9,
32'h3D282B97,
32'h3D66F3E9,
32'hBC3B9310,
32'hBD245F88,
32'h3D530DA3,
32'hBCBDB363,
32'h3D973BB7,
32'hBCF51341,
32'h0ECB581C,
32'hBDA83505,
32'hBD70891B,
32'h3DB0B015,
32'h3D25DFF8,
32'h3DCE6EE0,
32'h3C98A257,
32'hBC23CCD5,
32'hBA1A1CC,
32'hBD186E5A,
32'hBCB07135,
32'h3D839E07,
32'h3D770136,
32'h3C2A8A8A,
32'hBDA469B9,
32'h3D1187F5,
32'h3D9E5146,
32'hBD6882F1,
32'h3D2C1600,
32'hBDB3FC02,
32'h3D33E1E1,
32'h3C8150A1,
32'hBD8843B1,
32'h3D3890C5,
32'h3D3D9CCE,
32'h3D52432E,
32'hBC63C99C,
32'h5DE4BD18,
32'h3D03BB6A,
32'h3CFDA2D2,
32'hBC5A8786,
32'h3D71D034,
32'h3D00694D,
32'h3CB0C884,
32'hBD9C3154,
32'h3D89A0D3,
32'h3D273D71,
32'h3C14FD4C,
32'h3D5F8900,
32'hBC21C7B3,
32'hBC88F40E,
32'h3CB63772,
32'h3D0B4116,
32'h3D44D4E5,
32'h3D6A634D,
32'hBD03C020,
32'hBDD96144,
32'h3D9223AB,
32'h3DB418D6,
32'h3D5AE39E,
32'hBCDA0C6A,
32'hBC4C07B7,
32'hBCAB3614,
32'h3C14C438,
32'h3C8FFCC2,
32'hBD38E3CE,
32'h5DF5DC79,
32'hBCB6ED9E,
32'h5DD43BF2,
32'h3DAD81B3,
32'h3D9E5ACA,
32'h3D4C5860,
32'h3C8C6FDA,
32'h3D890D95,
32'h5DDCD466,
32'hBD02A3AB,
32'hBD010DBF,
32'h3CAE5A34,
32'hBCC23AB0,
32'h3C2E9B2A,
32'h3D929445,
32'h3DA2DD81,
32'h3D31A91E,
32'h3D14B71F,
32'h3D2EEB78,
32'hBD8C95D6,
32'h3C97ACFD,
32'h3D89A9D6,
32'hBC62DB39,
32'h3D577E93,
32'hBCB3D837,
32'h2E4ECC4,
32'hBD102F28,
32'h3CCE54F3,
32'h3DE9A9AC,
32'h3D0EF741,
32'hBCE2E454,
32'h3D5E83EE,
32'h1DF1A9CC,
32'hBC62CBED,
32'h0758DEB9,
32'hBDACE555,
32'hBC707538,
32'h3C8684C8,
32'h3D486885,
32'hBD3F6594,
32'h3D50979C,
32'h3D12DB25,
32'hBD96E718,
32'h3D37DE34,
32'h3D1B2A3C,
32'hBD3756B6,
32'hBCADE987,
32'h3D575B5F,
32'hBDAF59D6,
32'h3D6E5C3E,
32'h3DCCEEE9,
32'h3CF4C267,
32'hBD4FE6FE,
32'hBD84DF8F,
32'h3CB9D9F2,
32'hBD2B34A4,
32'hBD4927A7,
32'hBC9D04C9,
32'h3C9A1578,
32'h2ECE7669,
32'h1DC4716C,
32'h3C93D565,
32'hBC9ED878,
32'h3D074571,
32'hBDB259C4,
32'hBD0856FD,
32'h5DF505B4,
32'hBC6C65F8,
32'hBD228510,
32'h3C14E635,
32'h3D4EBCF0,
32'hBC0DDF21,
32'hBCF5F551,
32'h3C1D93F6,
32'h3DB56678,
32'h5DFC8CF7,
32'hBDDA5BCB,
32'h3D7EC61C,
32'hBD089994,
32'hBDA7ECEA,
32'hBCB00954,
32'hBC8ABD6D,
32'hBD8B2C3A,
32'h3D1C321C,
32'h3D02AC2A,
32'h3D936A8C,
32'h3C962A05,
32'h3D139DDB,
32'hBCC3BA55,
32'hBD0F4E59,
32'hBD2D1C6F,
32'hBDAEC6A1,
32'h5DFB6FF4,
32'hBC056B16,
32'h3DD99A25,
32'hBD8E9E05,
32'hBDB57A76,
32'h2EC743CF,
32'h3C94355A,
32'hBDAB8C4F,
32'h2ED7615A,
32'h3D468167,
32'h3D8BFF50,
32'h3D29377D,
32'h3A6B193,
32'h3D8A48C5,
32'hBCBED7FE,
32'h07595A21,
32'hBD67B716,
32'h3E275057,
32'h3CFB2F36,
32'hBCEF304E,
32'h3CBAE6E1,
32'hBD1BF540,
32'h3DA7B869,
32'hBD6BFF55,
32'h3D860259,
32'hBDFE10D5,
32'h3CC00AFD,
32'hBE1A0316,
32'h3D7EAEBF,
32'h3CBB14D9,
32'h3E1B11CD,
32'h3CCC0FA8,
32'h0ED06318,
32'hBD8B9EA8,
32'h3DB2D915,
32'hBD3B25ED,
32'h3CA7C815,
32'h3C6DEFDE,
32'hBDA92315,
32'h3C706F6B,
32'h3D86C093,
32'h3A0EF35,
32'h3D6AA13A,
32'hBD43E053,
32'hBC03BE84,
32'h3DB6A4A3,
32'h1DDD42FE,
32'h3DFAA419,
32'h3E1A8EA4,
32'hBE51FBC8,
32'hBD615CD9,
32'h3C75064F,
32'h3CDB2C20,
32'h3CEB540B,
32'h3CA8D5AE,
32'hBE291810,
32'h3D2DAE13,
32'hBE856ACA,
32'h3E68CD9A,
32'h3D04BCE8,
32'h3E3B32C1,
32'hBDA143F6,
32'h3E3BB1EE,
32'hBDCDEF4A,
32'hBCD019CA,
32'hBCD6382F,
32'hBC11E363,
32'h3C049BA5,
32'hBDB00C1E,
32'h3CFC887F,
32'hBD831F76,
32'h3D38F79D,
32'h3E21A882,
32'h3D4BBB17,
32'h3D223879,
32'h3DE13F23,
32'h1CEAE63,
32'h3E153FCE,
32'h3E6621B5,
32'hBE147444,
32'h3C959078,
32'hBD554D43,
32'hBD288D1E,
32'hBC6D44EB,
32'hBDCB874B,
32'hBE1ED1C5,
32'hBD926626,
32'hBE6CFB2A,
32'h3E5D2403,
32'hBDB04840,
32'h3E33CA15,
32'hBD0BE0D4,
32'h3CE0E0A1,
32'hBC914540,
32'h3D530DAC,
32'hBDA1E32C,
32'hBC11BA56,
32'h3CDA6CF6,
32'h3D00E169,
32'h3D091F4F,
32'hBD82C82E,
32'h3D2F4804,
32'h3DEAD0F4,
32'hBD5AFFBB,
32'hBC8EF8B4,
32'h3D7B212B,
32'hBCBE5BA8,
32'h3DE76E04,
32'h3C288896,
32'hBD55E055,
32'h3D7AF44D,
32'h3C875AC4,
32'h3D9E8A51,
32'h3DE0C319,
32'hBCC30055,
32'hBDA7DB04,
32'h3D845F23,
32'hBE2BCE63,
32'h1DC10F38,
32'h3CBA27E9,
32'h3D68802D,
32'h3D9C27CF,
32'h1DEC8C4B,
32'hBD20A49E,
32'h3C7966EA,
32'hBD45AC45,
32'hBD97AAF3,
32'hBDCE106B,
32'h3C827E56,
32'hBD968324,
32'h3C552136,
32'h3D727958,
32'h3C3F4383,
32'hBD96C57F,
32'hBCECEFFE,
32'h3DB7852E,
32'hBC9E84DF,
32'h3DCDA38C,
32'h3D460B34,
32'h3D9C867F,
32'h3DDE16BC,
32'h3C6A4054,
32'h3D59425B,
32'h3D32FEDD,
32'h3CE63EBF,
32'h3D013239,
32'h3D6DFDA4,
32'h3D138CEB,
32'h3CFB30E8,
32'hBD89A3DD,
32'h1DFD7F57,
32'h3D6DDDE3,
32'hBCD5F923,
32'hBC83DBDD,
32'h3CDEEDAE,
32'hBD8B4FB5,
32'hBCA65C99,
32'h3C6936CA,
32'h5DFE74CE,
32'h3C7B3DE0,
32'hBD5592B2,
32'h5DDDED26,
32'hBCBBCB4E,
32'h3CC9ED9B,
32'hBC14B3C7,
32'h3CDB1E96,
32'h5DD738AC,
32'h3D43107F,
32'h3DE8B3E3,
32'h3C0C0E95,
32'h3CAFEAF4,
32'hBDBD1566,
32'h0EC8D0AC,
32'hBDBEB34A,
32'hBD62E92D,
32'hBCAF1658,
32'hBCB8E371,
32'hBD1FECE5,
32'hBD3B75B1,
32'h3CFA04C6,
32'hBD156310,
32'hBCBDA790,
32'hBD26E8D6,
32'hBCBE0C73,
32'hBCFA516A,
32'hBCA40DB2,
32'hBCC5F040,
32'h3D4EFEB1,
32'hBCF49742,
32'h0EC570DD,
32'hBD8DEF06,
32'h3C3FB94F,
32'hBD8D3125,
32'h2ED6BA99,
32'h3D5F1452,
32'hBDBB64E5,
32'hBD30EDCF,
32'hBD62748F,
32'h3D368524,
32'h3D00BFA1,
32'h3D5F6AD1,
32'hBC27A076,
32'h3D8E39D0,
32'hBC5B9873,
32'h3CB60D35,
32'hBDC016AD,
32'h5DC37B68,
32'hBD0472D2,
32'h3C19C924,
32'hBD497AF8,
32'hBD4E34AA,
32'hBD71B6CF,
32'h2EDB2B76,
32'hBC503BAA,
32'h1DEA69A4,
32'h2EC97C70,
32'h3C260B03,
32'h3D9A26DB,
32'h3C8A6683,
32'hBD86D099,
32'hBD99153E,
32'hBD565DAF,
32'hBD671F81,
32'h3D647E45,
32'hBD44AFCF,
32'hBD11D7F6,
32'h2EC9C5D6,
32'hBD917920,
32'hBC9BC2EC,
32'h5DFEEB27,
32'h3C8F2831,
32'h3DBA300C,
32'h3D9D49CA,
32'h3D6666FF,
32'hBD252948,
32'hBDACC1FE,
32'h3D323CA7,
32'h5DDCD9C7,
32'hBD27649A,
32'h3D8F757B,
32'hBD46E2D0,
32'h3DAD2ADF,
32'hBD1A0142,
32'hBDB4D6DA,
32'h3D115267,
32'h3C65C81C,
32'h3C8CAB5F,
32'hBD4FF9AF,
32'h3DCC21C8,
32'h0ED70063,
32'hBD21A54A,
32'h3D4F224A,
32'hBD013EE2,
32'hBCDA853F,
32'hBD21D42B,
32'hBA48572,
32'hBDD95682,
32'h3D32907B,
32'hBD984F67,
32'h3CEAFD61,
32'hBC9FC67B,
32'h1DF14A78,
32'h3D268A38,
32'hBD78280A,
32'h3D19CC31,
32'h3C4FEC95,
32'h3D1127BE,
32'hBD5E4D54,
32'hBDBCABC6,
32'h3C4BBAB8,
32'h3DCE0030,
32'h0750BE0F,
32'hBC8D4BCD,
32'h3D0A1531,
32'h5DC3DA49,
32'h3D96B0AD,
32'h3C64B66E,
32'h3D4A52CB,
32'h3CAF26A7,
32'hBDD891D6,
32'hBCCB777B,
32'h3CD826F6,
32'hBD85DD54,
32'h3DC30775,
32'hBD29CBB4,
32'hBC80B6F7,
32'hBD9816B1,
32'h3D86303D,
32'hBD31CAFC,
32'h3C0F8313,
32'h1DFAB747,
32'h3CEB6A68,
32'h3C54EB65,
32'h3D69B9B2,
32'h3D643107,
32'h3CE5B55E,
32'h3D4E51DD,
32'hBCBDA9F5,
32'hBCB4D4BC,
32'h3C4DA177,
32'hBD0FB7C2,
32'h3D4D0704,
32'hBD699243,
32'h3D0D2868,
32'hBD344717,
32'hBCEA6EEC,
32'h1DEDABA5,
32'hBC64863D,
32'h2ED3156D,
32'hBCAB6873,
32'h3CB0883E,
32'h3C00A28F,
32'h3CFF8DCC,
32'h5DF5BC3C,
32'h3CB51745,
32'hBCCD4070,
32'hBD7A6853,
32'hBDD31AEA,
32'h5DF7BB86,
32'h3D4D8B50,
32'h1DC63A38,
32'hBDC01C6E,
32'hBD36E64C,
32'h3D2288A6,
32'h3D353345,
32'h3DC40D7C,
32'h3C24918E,
32'hBD4BA5B4,
32'h3DDE09B7,
32'hBC5BC926,
32'hBCEBE371,
32'hBC861B81,
32'hBD9923DF,
32'h3D9E2618,
32'hBC8E8FCE,
32'h3A6C0E6,
32'h3D263A58,
32'h175A079F,
32'h3C888F48,
32'hBD02BBBB,
32'hBD6F8E24,
32'hBD3BA317,
32'h3D9170AC,
32'h3C962DB6,
32'h1752825B,
32'h3C8B80A7,
32'h3C85FAB9,
32'h3D7BC6CB,
32'hBD25A3E1,
32'h3D203F06,
32'h5DEA4954,
32'h3D7DDEB8,
32'h3DA597D5,
32'h3D3CA7CA,
32'hBDA535E9,
32'h3D3F9DEE,
32'hBCB142EB,
32'h3DC21533,
32'h3D114F7D,
32'hBD051384,
32'h3CAE3A88,
32'h3D7F2B91,
32'hBCA5449F,
32'h3CAFCE80,
32'hBCF21D4E,
32'h3DCC28BD,
32'h3DB6BFA6,
32'h1DFA1A4E,
32'h3D002AD5,
32'hBC5DB306,
32'h17567AC7,
32'hBC699B55,
32'h3D237EAF,
32'hBCF2CA42,
32'h3D46420D,
32'hBD668A30,
32'hBD1FF62A,
32'h2EDBC343,
32'h3D39561C,
32'hBD170854,
32'hBD500703,
32'h3DCD6BEB,
32'h3C7DFDBA,
32'hBCB6FFC7,
32'hBC34D51B,
32'hBC0025E4,
32'hBC544719,
32'hBD9B3686,
32'h3C9D10E7,
32'h0757B2AD,
32'hBC05FD0E,
32'hBC943AEF,
32'h3C319A7C,
32'h3CCB560E,
32'h3CA014D8,
32'h3D81A7F0,
32'h3C1B04BC,
32'hBC6BC8A4,
32'hBD23566F,
32'hBDD26DEA,
32'hBC0F940B,
32'hBC775925,
32'h3DA99614,
32'hBD3174F7,
32'h3D75A583,
32'hBD86926C,
32'h3C7FA14D,
32'hBD186B3F,
32'h3D1D0ECF,
32'h3D0B4618,
32'h3D20E89D,
32'hBD994897,
32'hBC718456,
32'h3C34CA03,
32'h3CC68697,
32'hBD02F393,
32'hBCA97A02,
32'hBD9A527A,
32'h3D0F4D53,
32'h3DD803C5,
32'hBD947719,
32'hBD52FE16,
32'hBDC9DD5A,
32'h3CB9A14A,
32'h3DAABC99,
32'h3CD0E759,
32'hBC508D75,
32'hBC277DEF,
32'h1DFA3A2C,
32'h5DCFE74C,
32'hBD61DDBA,
32'h3D2EEFAC,
32'hBC18D627,
32'h3C89A2DC,
32'h3CB1BC89,
32'h3CDF828D,
32'h3D6A5048,
32'h3D215418,
32'h3DA5D48D,
32'hBC796F35,
32'h3DBD28BD,
32'h1DEC025C,
32'h2EDD577E,
32'h3D8CA12B,
32'h175249B5,
32'hBD22B249,
32'hBD7594FD,
32'hBC394124,
32'hBD2ED32A,
32'h3D7F0063,
32'hBD170AD0,
32'h3D77BDC1,
32'hBDAF259A,
32'hBDD99341,
32'hBD23B33F,
32'h3D3E20E1,
32'hBD816ADA,
32'h0756CFE5,
32'h3D3F5DF8,
32'h3C439A1D,
32'h3CBD899C,
32'hBCB04B72,
32'hBCAD2DD0,
32'hBD3FD60C,
32'hBD03F957,
32'h3D8083C3,
32'hBD1023BF,
32'h3D93C925,
32'h3D3F077D,
32'hBCCEB515,
32'hBDAC33F4,
32'hBD13D20F,
32'hBC8EE2F0,
32'hBCA33573,
32'hBDBEFA28,
32'hBD7267FC,
32'hBD171FFB,
32'hBCD21C8A,
32'hBD57F0C3,
32'hBD54E136,
32'hBD44E526,
32'h2EDD0639,
32'hBDDC9871,
32'hBD07C8F1,
32'h3D217481,
32'h3D5CB472,
32'hBC34FB82,
32'h3D516050,
32'h3D61C33B,
32'h3DBE4258,
32'h3D8533A7,
32'hBDB237FB,
32'h2E58DF7,
32'hBD7239A0,
32'h3D6174D3,
32'h3D3BCD6C,
32'hBCBEA41D,
32'hBD5FED8C,
32'hBD2B4C5F,
32'hBCF76D57,
32'h0ECCF2BA,
32'h3C0CB333,
32'h3D205360,
32'hBCBEC5BB,
32'h3CB70A3B,
32'h3CDB1E2B,
32'h3DDB88D9,
32'h3D65091B,
32'h3DC478E0,
32'h3D29382A,
32'hBD0815FC,
32'h3C6D5BF7,
32'h3DAF695C,
32'hBC825300,
32'h3DA4CE28,
32'hBCC71F3E,
32'hBD2341FB,
32'h1CCA032,
32'hBC7C05B5,
32'hBC59C42C,
32'hBC1B6B7F,
32'h3D877475,
32'h3DB1EB3F,
32'hBDB6696D,
32'h3D25F87A,
32'h3DA68BC6,
32'h3D75A890,
32'h3CD8E1D3,
32'h3D201736,
32'h3D218B39,
32'hBCDBC661,
32'hBDBF0CC1,
32'hBCF81041,
32'hBD65059C,
32'h3D1998BD,
32'h3D35F5EF,
32'h3DC4AECA,
32'h3D11384B,
32'hBD377A0C,
32'h5DE79F06,
32'hBCBCCA83,
32'h3D401625,
32'hBD234366,
32'h3C8D24DE,
32'h3CA20145,
32'hBCAE0AC3,
32'h3D3085A4,
32'hBCA36FC1,
32'hBD8A80B9,
32'h3D98E0A9,
32'hBC8B5E83,
32'h3C0D1FB3,
32'h5DCC502E,
32'h3C8FC03A,
32'h3D23F38A,
32'hBD2399A8,
32'h3D317E56,
32'hBCEF6888,
32'h3C6A5FEF,
32'hBC313F25,
32'hBCD9059E,
32'h3C676B90,
32'h3D3A58F7,
32'hBCB9323A,
32'h0ECF4AB7,
32'hBDC77C16,
32'hBCB2128D,
32'h3A690BB,
32'h3D167395,
32'h3CF3B862,
32'h3DA3E146,
32'h3D3038E7,
32'h3C1F4F60,
32'h3DE7976B,
32'h3C8894EF,
32'h2ED8391C,
32'h3DACF5F2,
32'h3CDAE3C2,
32'h3C88277F,
32'h3D1C006C,
32'hBDB68AE6,
32'h3D45D698,
32'hBD50E14E,
32'hBD5C3961,
32'h2ECBFDE4,
32'h3D273901,
32'h3C73552E,
32'hBDE47016,
32'hBD8541A1,
32'hBD3410C0,
32'h3C8F633F,
32'h3DAE81B0,
32'h3C7D68A3,
32'hBCAC29EA,
32'hBCC0F763,
32'h3C9797DF,
32'hBDCDEB50,
32'h5DC45673,
32'h3C9A533D,
32'h5DE6CC5D,
32'h3D77415D,
32'h3D118940,
32'h3D45C951,
32'h3DCB3288,
32'hBD2A8866,
32'h3D4869D6,
32'hBDB3168C,
32'h3C89EA44,
32'hBDE42E5B,
32'h3DA6D07D,
32'hBD79B8E6,
32'hBCC1C891,
32'hBCDC17C1,
32'h3D539EDE,
32'h5DE11CCE,
32'hBD3512C2,
32'h3CDA5726,
32'h3C8842A6,
32'h3D2B53DF,
32'hBCDA2613,
32'h2EC05AAD,
32'hBD8A0DDD,
32'hBCC7E027,
32'hBD07DCA9,
32'hBC559915,
32'h3D4BCB99,
32'hBD268B06,
32'h3D4C5391,
32'h3DDD3DDF,
32'h075AFA45,
32'hBCFEAFDD,
32'hBC06399A,
32'h3D40AC6D,
32'h3CD0E2BB,
32'hBC853210,
32'hBD983F76,
32'hBD496B40,
32'h3D502F0E,
32'h3D91AF6A,
32'h3D7833EC,
32'h3CD2182A,
32'hBD552AD2,
32'hBC76A329,
32'h3C44D04C,
32'h3CC7B9DE,
32'h3D45C0B1,
32'h3DEFAC0E,
32'h3C97E13A,
32'hBDAECA1A,
32'hBDBE56AD,
32'h2ED93879,
32'h5DDCBF99,
32'h3CFFF37F,
32'hBD6D8A12,
32'h3D1D490E,
32'h3DC3F3B1,
32'h3D0139C6,
32'h3D8F4FF8,
32'hBDE7273B,
32'h1DC97FE1,
32'h3D804F8E,
32'h3D76FD95,
32'hBD3EFBF2,
32'hBDF28AE2,
32'hBD339291,
32'h2ED284AE,
32'h3D4EAE7D,
32'hBD50A4FA,
32'hBD13BF60,
32'hBDD830E5,
32'hBE0A80D5,
32'h3D37A053,
32'hBE807117,
32'h3C7DAC56,
32'h0EDF7CCA,
32'hBD4B3EAF,
32'h3E690308,
32'hBC83A366,
32'hBD3FFD54,
32'h3D869650,
32'hBD90CF04,
32'hBD80D068,
32'hBE6318CB,
32'hBECB32A2,
32'hBDC2ACC7,
32'h3EFC807E,
32'hBD95ADC5,
32'h3ECB6EA9,
32'hBDC9C41F,
32'hBE252C94,
32'h3E6FA464,
32'h3D9A8A4F,
32'hBD9EE856,
32'hBE5EBEF7,
32'h3D89CE9C,
32'h3C753FB1,
32'h3A37773,
32'hBCBB8528,
32'hBD8B8CE5,
32'hBCB314E3,
32'hBD2D64A3,
32'h3CCEA803,
32'hBEA4D45B,
32'h3A02F7E,
32'hBDCC5C86,
32'hBD72C337,
32'h3E93C1C6,
32'hBC8C6C97,
32'h3D436E15,
32'h1DDB50AE,
32'h3E00566F,
32'hBDF9D67E,
32'hBE8CA517,
32'hBEC52903,
32'hBE1E7ABD,
32'h3EADFF9C,
32'h3D5BA476,
32'h3EF860F6,
32'hBDAD7DB6,
32'hBCA7FC55,
32'h3C896659,
32'h3D0EC077,
32'hBE78C042,
32'hBE272293,
32'h3DAFAB17,
32'hBD399399,
32'hBD5551EE,
32'h3E17DDA8,
32'hBEA6BDDE,
32'h3D715739,
32'hBEE97BF3,
32'h3DFF22A2,
32'hBDF2253A,
32'hBA438CE,
32'hBD15004D,
32'hBCAF0EB4,
32'h3F15F7A6,
32'hBDEE0490,
32'h3CB76C84,
32'hBD8BC901,
32'h3D8A6304,
32'hBDCE70CB,
32'hBDE2CBFC,
32'hBE7C8D92,
32'hBDE426DA,
32'hBC85B306,
32'hBE220D88,
32'h3F35A1BA,
32'hBDD03F8A,
32'hBD0324FF,
32'hBE4627BE,
32'h3CE2EA3D,
32'hBDB0242F,
32'hBDC63419,
32'h3D0FE1ED,
32'hBD1E7C80,
32'hBC6FD95B,
32'h3F5A6DDA,
32'hBEF100DD,
32'h3D6D8A06,
32'hBFAAB745,
32'h3DB3EA4A,
32'hBEBA5F3C,
32'hBDE19543,
32'hBC8F83DC,
32'h3CCB6437,
32'h3ECED806,
32'hBFB29731,
32'hBD942F36,
32'h3F24991E,
32'h3DCFA2B5,
32'hBE6011DC,
32'h3D7AC762,
32'h3EDB0C1F,
32'hBD5406A4,
32'h3E5714BB,
32'hBE1D0C96,
32'h3FADFE01,
32'hBEA49B83,
32'hBDE9330A,
32'h3E635E57,
32'hBD6FBBC6,
32'hBF3B98A0,
32'h3DB447A9,
32'hBD02797A,
32'hBD10E100,
32'h3F203210,
32'h3F665AC9,
32'hBE2B1E3B,
32'h3CC06A2B,
32'hBF424982,
32'h3ECF796B,
32'hBF094C1C,
32'h3C6C0AD1,
32'hBD927697,
32'h3D39C5C4,
32'h3E53ABE6,
32'hBF7D7D67,
32'h3EFEB871,
32'h3F234AD3,
32'h3E05C132,
32'hBE621247,
32'h3D9B2162,
32'h3EFD45AA,
32'hBD932696,
32'h3DB56078,
32'hBD379224,
32'h3FB825FC,
32'h3E2F7F09,
32'hBD723F6D,
32'h3F1AA587,
32'h3C9BFF53,
32'hBF235591,
32'hBDE1EE53,
32'hBC7D4180,
32'hBD07B964,
32'h3EC5A599,
32'h3E569601,
32'hBE8C911E,
32'hBEA26887,
32'hBCD5BEC8,
32'h3FBB0FD2,
32'hBDFF3C61,
32'hBF04DBF9,
32'h3A5DC0B,
32'h3D41F535,
32'h3FC1A3BD,
32'hBEDA661C,
32'h3F24FB63,
32'hBF98EFAF,
32'h0EC372E5,
32'hBF3B4BE2,
32'hBE3B7893,
32'hBF824C0D,
32'hBF500F89,
32'hBD9F5758,
32'h3F789205,
32'h3F2F238B,
32'h3E96B71F,
32'hBCDBF473,
32'h3F8B1A94,
32'hBC263A56,
32'h3C722E08,
32'hBE9FB3B6,
32'hBCFE8B46,
32'h3A2AF7E,
32'h3E4447A2,
32'hBD2F63E9,
32'hBD192863,
32'hBE86DF1D,
32'hBE6E31BE,
32'h3F647B6E,
32'hBE3DD2EB,
32'hBEA03808,
32'h3C693163,
32'hBD812780,
32'h3ECA5A1F,
32'h3D526705,
32'h3F12BC8A,
32'hBF1225F4,
32'hBD002064,
32'hBE9FD82C,
32'hBD2430CE,
32'hBD9C0A98,
32'h3CFED3F9,
32'h3D8FF667,
32'h3F5065E6,
32'h3EF67F43,
32'hBE17C9C4,
32'hBD4613AF,
32'h3E0134AE,
32'hBD39FB5C,
32'hBE3FAD7C,
32'h3E85B4B3,
32'h3D169424,
32'hBCE0ADC7,
32'hBE62DDC9,
32'h3E087CEE,
32'hBD8E4F7A,
32'hBF063DD1,
32'h3F204B5C,
32'h3FDC0A22,
32'hBE1EB693,
32'h3EA618A0,
32'h3D06B77F,
32'hBCD0E3F2,
32'h3F2C5ADC,
32'hBE142D0A,
32'h3E6C5D3D,
32'hBEB74F51,
32'h3FA1ACEE,
32'hBF7D1C54,
32'hBF23313E,
32'h3E488DDD,
32'hBEDA2984,
32'hBE808795,
32'h3E80D598,
32'h3EF2D9AD,
32'h3CB58443,
32'hBD140EF8,
32'h3F0A052D,
32'hBDA3A31C,
32'h3F5BDAC9,
32'hBDA07E17,
32'hBE3B4373,
32'hBDF9097C,
32'hBE948B43,
32'h3E49CEF8,
32'hBD5989A0,
32'hBE068329,
32'hBE7B3A13,
32'hBE90F5FA,
32'hBCF97785,
32'h3E82318D,
32'hBCAEDBC0,
32'h3DC71E63,
32'h3E7F124D,
32'hBEEEBB93,
32'hBE268E87,
32'hBDF4DF20,
32'h3F929F64,
32'hBDFFB5BC,
32'hBE75317A,
32'hBE63B306,
32'hBCC1EB7A,
32'hBE3BD6A0,
32'hBEF8EEE8,
32'h3F2C28C8,
32'hBDDB38E1,
32'h3CC444AC,
32'hBE6DFED9,
32'hBD7E5178,
32'hBD5F1B8F,
32'h3F175E07,
32'hBEC1EE4B,
32'hBE8A3000,
32'h3E029DF0,
32'h3D3D9E0C,
32'hBE5BB66C,
32'h3CC79BCF,
32'hBEC8C766,
32'hBF0B5B43,
32'h3EB801DE,
32'hBE22FEB6,
32'h3C90C3D5,
32'hBCB501A1,
32'h3F3D56E0,
32'hBE649E49,
32'h3E7DFBE8,
32'hBF031D97,
32'h3FBDF509,
32'hBF81AD7F,
32'hBFC836C4,
32'hBFA49672,
32'hBEB29EEE,
32'h3E264118,
32'hBE8600AF,
32'h3F92EE8B,
32'h3D521D67,
32'hBEA9F242,
32'h3C872D6B,
32'h3D76E0BF,
32'h3E1B89E6,
32'h3F0A03FD,
32'hBFC5A451,
32'hBDD576FA,
32'h3FA301BA,
32'h3E4BE5FC,
32'h3DFDDE95,
32'h3D3C7B85,
32'hBF07945A,
32'hBE41AEFE,
32'h3F8D6130,
32'hBF78FDD3,
32'hBC6B4BA8,
32'h3C4CB29A,
32'h3EF3FE41,
32'h3F146510,
32'h3FB5837C,
32'hBF91EF7E,
32'h3F7EE21C,
32'hBD91ADEF,
32'hBF5D750D,
32'hBF9913CF,
32'hBEB44575,
32'h3E9FAB9E,
32'hBF9B5F44,
32'h3EC728ED,
32'h3F2681D0,
32'h3D82FDA4,
32'h3E283F85,
32'h3D4A8080,
32'h3F86423E,
32'hBE5AF2F8,
32'hBE972FB9,
32'hBCF44296,
32'h3F642F92,
32'h3E52E8C2,
32'h3E80530D,
32'h3E2282DF,
32'hBE1E8525,
32'h3E893165,
32'h3DE96F30,
32'hBE111253,
32'hBDC24E07,
32'hBDA1DF5A,
32'h3F7A37E5,
32'hBC5873D2,
32'h3EBF1E29,
32'hBF544356,
32'h3F629F27,
32'hBDC8B186,
32'hBD989AC7,
32'hBF8A5B76,
32'hBE5B08CE,
32'h3E002A89,
32'h3EA665EA,
32'h3ECFA7E8,
32'hBE26C362,
32'h5DF9774E,
32'h3E0FC58C,
32'h1DC566A0,
32'hBE67D6E7,
32'h3E03807A,
32'h3D831C95,
32'h3C04ACCF,
32'h3E379753,
32'hBEA3F7FF,
32'hBD8D32AE,
32'h3D2326E2,
32'hBD90FCBE,
32'h3E8E7AE8,
32'hBE550C12,
32'hBF36B2CE,
32'hBD091962,
32'h5CC3C62,
32'h3F902441,
32'hBE14D20C,
32'hBE322205,
32'hBFDABE2C,
32'h3EF9BFB3,
32'h3DCC9DFB,
32'h3DDF8D2C,
32'hBF0E2C72,
32'hBE7E159A,
32'hBEAFFD91,
32'h3F94C701,
32'h3F09E808,
32'hBDC1932B,
32'hBD7D0F9A,
32'hBEEFC6C7,
32'h3F52C0B1,
32'hBE63F5AE,
32'hBCEE0475,
32'h3D5C0E68,
32'hBC54418D,
32'h3CBB47FB,
32'h3D9C438D,
32'h3D2BCC3D,
32'h3E869703,
32'hBEEF4E2A,
32'hBE42202A,
32'h3F1E48F1,
32'h3D026092,
32'h3DCF621C,
32'hBD223D72,
32'h3F5696A9,
32'h3D42C83B,
32'h3D9CF060,
32'hBDDE3C17,
32'hBD4572CE,
32'h3CEF5F70,
32'hBF0F5A12,
32'h3EE9D314,
32'hBDCE1DAC,
32'hBE0C2246,
32'hBE91974C,
32'h075153FA,
32'h3D0ACC94,
32'h3D7B766D,
32'hBDBC2E36,
32'h3D2D8E48,
32'hBDA75C35,
32'h3DE67525,
32'hBC9E1E14,
32'hBC3AC621,
32'h3C235D1C,
32'h3C685A7D,
32'hBC8857C0,
32'h3EA06C7D,
32'hBD9A396E,
32'hBDF21E70,
32'h3F0B03B6,
32'hBD130B3F,
32'h3E11B381,
32'hBD441B70,
32'h3F534EEF,
32'h3C4C380C,
32'hBD99004A,
32'hBE8E95AD,
32'hBCE296D3,
32'hBDE7D826,
32'hBECA74FB,
32'hBED3DC13,
32'hBE4ED6F1,
32'h3D3C3701,
32'h3ECD9B2D,
32'h3E87FAEB,
32'h07521A52,
32'hBD2CD00F,
32'h3D51D9A1,
32'hBD6E4749,
32'hBD62398A,
32'h2EC623DF,
32'h3DA43021,
32'h3DB11107,
32'hBC22C542,
32'hBC14E9DE,
32'hBCE738F9,
32'h3EE50434,
32'hBECA336B,
32'hBE4B48B2,
32'hBD97D138,
32'h3C0F2E84,
32'h3CEF3CE7,
32'hBC13C2F7,
32'h3F276D54,
32'hBE283F7B,
32'hBE40544B,
32'hBC8C8AC9,
32'h3D6F987D,
32'hBD9EB86C,
32'hBE41D094,
32'h3E138C36,
32'hBD5B0F6B,
32'h3E0575B3,
32'h3E40D755,
32'h3D1BA13E,
32'h3DECCC60,
32'hBA2748A,
32'hBE401661,
32'h3CB38DC0,
32'hBC5AB015,
32'hBCE1E069,
32'h3D84CFDD,
32'h3D194051,
32'h3DC670F5,
32'h5DDA727A,
32'hBE0AB35E,
32'h3EC9F361,
32'hBE8B46C4,
32'hBEC78F00,
32'hBE79B9F8,
32'h3E015955,
32'h3D99EEF5,
32'hBDDB0D26,
32'h3F617290,
32'h3D0ABA35,
32'hBE426C60,
32'h3D41A357,
32'h3D88B835,
32'hBD06B80B,
32'hBE8F9CE7,
32'h3E729CE0,
32'hBDBF72F1,
32'h3D04CAC2,
32'h3DED1EB6,
32'h3E2E74BB,
32'h3E8AD846,
32'hBD0D1597,
32'hBE4697ED,
32'hBDA2AED2,
32'hBD47BEBF,
32'hBE3BA611,
32'hBD5FC76D,
32'h3D6FB2C4,
32'h5DC87E2F,
32'h3D9B87CB,
32'h3CC8F19E,
32'hBD938372,
32'hBD15DD60,
32'h3CE0DED5,
32'hBD862FA2,
32'hBC89D264,
32'hBDE36F48,
32'h3D106E7D,
32'h3E07D0EF,
32'hBD4E663B,
32'h3D184338,
32'hBD9B01DC,
32'h3CC1E374,
32'hBDEDD5FA,
32'hBDC86F74,
32'hBD0F3EA9,
32'hBE17B54A,
32'h3DD163E5,
32'hBCDF5700,
32'h3D0F00BC,
32'h3C802CC5,
32'h3C908496,
32'h3D3D8EED,
32'h5DE2435B,
32'hBCC7F6B3,
32'hBD3439BF,
32'hBD464D6E,
32'h1DD1016A,
32'h3DC11770,
32'h3D81E009,
32'hBC47072A,
32'h3C95D909,
32'h3C609C07,
32'h3D1D14F5,
32'hBC9D51A2,
32'h3D805156,
32'h3DC46D08,
32'hBD3C8719,
32'hBD7C49DB,
32'hBC2CAB23,
32'hBDB66CF7,
32'hBD44F892,
32'hBCC4B4E3,
32'h3D263D3B,
32'h3C1C39A7,
32'h3C94BAAC,
32'h3C9FC499,
32'hBCC0A731,
32'h3D6C1AE6,
32'hBD8B2D32,
32'h2EC14F20,
32'h3C7BF5D2,
32'h3D7ABD38,
32'hBDB8A69A,
32'hBC959660,
32'hBD8868BE,
32'h3CB3C49F,
32'h3CDC4F18,
32'h3D78B110,
32'h3CD6C1E8,
32'hBD2F4B5D,
32'hBD06E9B9,
32'hBC74EE71,
32'hBD8A5E81,
32'h3CFFF487,
32'h3D56F590,
32'h3DD95AC0,
32'h3CD72605,
32'h3D249554,
32'h3C57D850,
32'hBD02F9BE,
32'h3D16F4E1,
32'hBDE9AFF5,
32'h3D9733FA,
32'h3D967E70,
32'hBD5A2A51,
32'h3C90BEBC,
32'hBCB50BF0,
32'h5DD44EA0,
32'hBCC2EB09,
32'hBDBC693B,
32'hBC1E9C44,
32'h3CBB4405,
32'h3DA2C262,
32'hBD17B4BB,
32'hBD3422E5,
32'h3D151894,
32'h3D89F7DD,
32'h3DC68861,
32'h3C74221E,
32'h3C5DF82B,
32'h3D2DE35A,
32'hBC5139B2,
32'h3D15342B,
32'hBDB8F14C,
32'hBD73A105,
32'hBD83238F,
32'hBCB5C580,
32'hBD97A97C,
32'hBCE9D2DC,
32'hBD8854CC,
32'hBCEF9450,
32'hBC41F6BD,
32'hBD048E47,
32'hBDC6561C,
32'h3DA2FAFD,
32'h5DF22C95,
32'h1DDB6EFC,
32'h3DB17856,
32'hBD4F7DC1,
32'h3DB076FF,
32'h3CA280B9,
32'h075D217D,
32'hBD061F37,
32'h3DA346BC,
32'h3D08C135,
32'h2ED673C7,
32'hBD07647F,
32'h3D2CF0EF,
32'hBA3C8E3,
32'h3CC74005,
32'h3D24A083,
32'hBA1CB26,
32'h3D3960C7,
32'hBD14B225,
32'hBD47584E,
32'h3DA72EF6,
32'hBC3D6AC9,
32'hBCE79520,
32'hBCE4307B,
32'h3D7F13BC,
32'h3CEE6FDA,
32'h5DF1A142,
32'hBD0E7999,
32'h5DCB569E,
32'h3D9C1275,
32'h5DEA7EBE,
32'hBCA12E59,
32'h3D5228AC,
32'hBCE862AE,
32'hBCA54C89,
32'h5DCE13D7,
32'hBCD563CA,
32'h3DA87712,
32'hBD739588,
32'h5DD019C3,
32'h3C866843,
32'h3DBC22CC,
32'hBD258A29,
32'hBD43F940,
32'hBD809EA2,
32'h3D70C2C0,
32'h0758F558,
32'hBD181FFE,
32'h3D2D1326,
32'h3D9A7C78,
32'hBC8204CF,
32'hBD5DCCF4,
32'h3D7A3042,
32'hBCDBC1C7,
32'hBC5B7959,
32'hBD191039,
32'hBD5CF464,
32'h3C4E7A60,
32'h0ECF6F05,
32'hBC10D58B,
32'hBDB8B862,
32'hBDE5F8E4,
32'h3CF76C6D,
32'h3D217ABC,
32'hBDE44274,
32'h3D1B8561,
32'h3D233523,
32'h3D90F9F4,
32'hBC613DB9,
32'hBD85729E,
32'hBC7CCC03,
32'hBD192367,
32'h3D047DFC,
32'h3C4948C8,
32'h3D7C6175,
32'hBD084CE0,
32'h3C4C787A,
32'h3C8E4A9F,
32'h3D6A131B,
32'h3DACC44F,
32'hBC6DAEC2,
32'hBD220DEF,
32'hBCF08F0E,
32'h3CFFD35B,
32'h3D30AA83,
32'h3D3DBA50,
32'h1DE83BC7,
32'hBD1FE665,
32'hBDB35900,
32'hBD8F0C0A,
32'h3DB75AE8,
32'hBD3064C0,
32'hBDAFD22D,
32'hBD512F33,
32'h5CC9179,
32'h0ECC5920,
32'hBD7B5A0D,
32'h3CDC0963,
32'hBD79B5AB,
32'hBCEAED86,
32'hBD8D87D5,
32'hBCBF434C,
32'h3C8F57D1,
32'h3D0AF598,
32'h5DF01DA9,
32'hBCCD33D0,
32'h3C9E6312,
32'h3D17CBE3,
32'hBCFE6308,
32'h3D98B785,
32'h3DBA9510,
32'h3C4411FA,
32'h3CE666F1,
32'h3CE4ABA1,
32'h3D964D88,
32'h075F3FFC,
32'h3CE3BF8E,
32'h5DC2A656,
32'hBD905661,
32'h3D91F96F,
32'hBDDEB4AB,
32'h3D5B455D,
32'hBD71732F,
32'hBD808650,
32'h0ED8348E,
32'hBCF5583E,
32'h3C1BC65D,
32'h3D0DCD15,
32'h3D43C752,
32'h3CDA0263,
32'hBDC6C5FA,
32'h3C16983E,
32'h0ED347FC,
32'h3EA2AEDF,
32'h3D173403,
32'hBDB3EEFC,
32'h3D19C02E,
32'h3E76E75D,
32'hBC1F3E6C,
32'hBCBD843C,
32'h3C8F19E8,
32'h3CF01B75,
32'h3ECF3F24,
32'h3D104291,
32'h3CC4CB74,
32'hBEA051A6,
32'hBCCF47FC,
32'hBD895CA1,
32'hBDF9F974,
32'hBEAC2CFB,
32'h3D86025C,
32'h3CDF3F70,
32'h3CCADB0D,
32'h3DBA3E05,
32'h3A2C784,
32'h3D8EBBDE,
32'h3D2BF604,
32'h1DE97EB2,
32'hBD221C33,
32'hBECBEACC,
32'h3C7883B9,
32'hBC937CFA,
32'h5DEABEC5,
32'h3E890735,
32'hBD211AA2,
32'h3DD93C0F,
32'h1DCAD372,
32'h3E522634,
32'hBCE59C77,
32'hBD324158,
32'hBCEFAE16,
32'h3CF8FA59,
32'h3EBAE96A,
32'hBC376965,
32'hBC7B7B3A,
32'hBEB7F063,
32'hBD42BC73,
32'h3C9335EA,
32'hBDED251D,
32'hBE7405DA,
32'hBC9E7EEE,
32'h3DE2946C,
32'hBC6A6B19,
32'h1DDE2745,
32'h3DAB5E07,
32'hBD907973,
32'h3D75C6C0,
32'h0ED3C1B4,
32'hBCABB71C,
32'hBEBAF6CF,
32'hBCE101E4,
32'hBD16E874,
32'h3DA4C9A0,
32'hBD8B30AB,
32'hBD9775C2,
32'h3D2AA77A,
32'hBD0DE78B,
32'hBDFF5B70,
32'hBDDA7093,
32'h1DE842ED,
32'hBD5B6388,
32'hBD06C58E,
32'h3E2CD14B,
32'h3E4B42C6,
32'h3DDC9D54,
32'hBD420067,
32'h3DF1D29C,
32'hBD28FDA7,
32'hBD758FCE,
32'hBE3B4BA4,
32'h3CC9F6B0,
32'h3DC8B567,
32'h3D3668F2,
32'hBD4A83BD,
32'h3E06E982,
32'hBDC80EC9,
32'h3E2CE6F2,
32'hBD32243C,
32'hBCB30C73,
32'hBE5CE313,
32'h3DBF9B15,
32'h3DDB4FB7,
32'h3EB37A9E,
32'hBDF7C278,
32'hBDC64B0B,
32'h3DB3B267,
32'hBD9E5829,
32'hBDE1E8BE,
32'hBD9C3FC6,
32'hBDC753E4,
32'hBD439800,
32'hBDC959E3,
32'h3E9E0350,
32'h3EB76922,
32'h3E0E65C8,
32'hBE3BF327,
32'h3E847489,
32'hBE30D792,
32'hBE601BB0,
32'hBE55C0A5,
32'hBD2450AC,
32'h3EA7203F,
32'hBDC1AC96,
32'h3F12B50E,
32'h3D460DB9,
32'hBD5A8674,
32'h3E1A7D71,
32'hBC898EFC,
32'hBE3744A1,
32'hBEC970B8,
32'h3D94A4AD,
32'h3E03D516,
32'h3E6E5EB0,
32'hBE94A8BD,
32'hBE2BF1F9,
32'h3D308A91,
32'h3EF04A4A,
32'h3F3C1E23,
32'hBE6503F3,
32'hBCCCB03A,
32'h3D2EC69E,
32'hBD0D0B57,
32'h3E3A6AFC,
32'h3F732F39,
32'h3EA0FA28,
32'hBCD30838,
32'h3ED17423,
32'hBDC29F8B,
32'hBE948CDB,
32'hBEBFC8E9,
32'hBDE65C39,
32'h3E98D7EA,
32'hBE799798,
32'h3F28CA07,
32'h3E01203C,
32'hBC87D80C,
32'hBA52484,
32'hBD3C2EAC,
32'h3E1EB135,
32'hBE950DCE,
32'hBCE06798,
32'h3CFD7477,
32'h3E7C29CB,
32'h3E7FB8F0,
32'hBF0B9A50,
32'hBF45EA22,
32'h3F291FC2,
32'h3EB22454,
32'h3E2E2403,
32'h3F50CF81,
32'h1756CDB0,
32'h3DD89532,
32'h3F53ABA7,
32'h3E09C341,
32'h3DB23521,
32'h5DEB41DF,
32'h3FE7AB0A,
32'hBE968C01,
32'hBE2C84D6,
32'h3D57D41B,
32'hBE2602AF,
32'hBEEFD3EE,
32'hBE88F1D7,
32'h3F42F8DD,
32'h3F243983,
32'hBDC60C0D,
32'hBE125D1C,
32'hBE69AF67,
32'h3E9CA806,
32'hBE37F019,
32'h2EC66A47,
32'hBE09CF29,
32'hBD665F6A,
32'hBFF25931,
32'h3EC4C645,
32'hBF15A0E2,
32'h3F3851E6,
32'hBE350975,
32'h3EF240A8,
32'h3E949E9D,
32'hBD114798,
32'h3D6FA2CA,
32'h3F9F2DD3,
32'h3ECE4E88,
32'h3EDF2F09,
32'hBF01B839,
32'h3FD22286,
32'hBE87FAE6,
32'hBE805B6E,
32'h3EC33D94,
32'hBE18B57B,
32'hBF0CF407,
32'hBF27F07E,
32'h3FEE8F9C,
32'h3E4512EF,
32'h5DC02787,
32'hBF100CAE,
32'hBEBA8F72,
32'h3F6B8261,
32'h3E6E7F6D,
32'h3DB75467,
32'hBE235DC2,
32'h3E649FB4,
32'hBE402C89,
32'hBF0DE109,
32'hBF7CDE25,
32'h3E3DC1FB,
32'h3F83F7E3,
32'h3D3D9C39,
32'h3F0CEA74,
32'hBDCC674F,
32'h3C7A40E9,
32'h3F99487D,
32'h5DFC76D7,
32'h3F3F86EA,
32'hBF2276DD,
32'h3F374197,
32'hBF06B05B,
32'hBF3009C3,
32'h3E78BC63,
32'hBF5CD049,
32'h3DB782FF,
32'hBEA22263,
32'h3FD30E98,
32'h3F12A27B,
32'hBD168AEE,
32'hBE6A5564,
32'hBE924031,
32'h3F8154FF,
32'h3ED7652D,
32'hBC9122C6,
32'hBEB311DD,
32'h3F29B8D0,
32'hBF62E24C,
32'hBE3F3FEF,
32'hBF0F0079,
32'h3F5EFDC3,
32'h3F6B66E1,
32'hBD90EB10,
32'h3F64A6D7,
32'hBD758D92,
32'hBD879329,
32'h3F6FA6DD,
32'hBD940B7A,
32'hBD327234,
32'hBF54D851,
32'h3DBCE68A,
32'hBFBE53B3,
32'hBFCC76A4,
32'h3E1E1845,
32'hBF69E105,
32'hBD4F8AD8,
32'h3E03F763,
32'h3FD0BC12,
32'h3ECA80AA,
32'hBE00CA95,
32'h3E85C730,
32'hBF139DB0,
32'h3F916C4F,
32'h3F3E67DC,
32'hBED0797A,
32'hBE2DE032,
32'h3FC42AB8,
32'h3CC56B14,
32'hBD5B72D3,
32'hBFCFBAD6,
32'h3E875BC5,
32'h3D67E7B4,
32'hBDFF4635,
32'h3E2A5F36,
32'hBDB2654D,
32'hBD3ABF0D,
32'h3FE64C3E,
32'hBE5A27FA,
32'h3D34DF95,
32'h3ECA607C,
32'h3EACC02F,
32'hBF8A13AB,
32'hBFD86F9F,
32'hBF0905D9,
32'hBF10B10B,
32'h3EC6D6B3,
32'hBFC3D526,
32'h402A8EE5,
32'hBECE661A,
32'hBD946F7D,
32'h3F77993B,
32'hBE58743D,
32'hBDD08954,
32'h3EFECE87,
32'hBEC56FA1,
32'hBEB9ED17,
32'h3EA3121F,
32'hBEE615E9,
32'hBE84A576,
32'h3E1CF80F,
32'h3E6BA460,
32'hBC831132,
32'h3DB245B5,
32'h3F627537,
32'h3D9B2E55,
32'hBDCB5E3F,
32'h3F7B3F14,
32'h3EA5D767,
32'h3EA10B76,
32'hBE83EC7A,
32'h3F95B71A,
32'hBF82CD27,
32'hBFD5E681,
32'hBF05CB49,
32'hBF1FAA0A,
32'h0EC97758,
32'hBFB04BB7,
32'h40025F61,
32'h3F01AD4B,
32'hBCFC529A,
32'h3D5216ED,
32'h0EC76A09,
32'h3F80C823,
32'h3F07EC2B,
32'hBEF71A17,
32'hBF4B8D79,
32'hBF266E2A,
32'hBFB4CB8B,
32'hBEADEF7E,
32'h3D9A6C44,
32'hBF1A03CC,
32'h3E269B5D,
32'hBF3831B5,
32'h3EB482F0,
32'hBD8893E0,
32'hBD05E164,
32'h3F07FBB5,
32'hBEB8FCE4,
32'h3F3920A0,
32'h3E066AE1,
32'h3E415C56,
32'hBFA1149C,
32'hBFD8864A,
32'h3F5FA696,
32'hBF9897BB,
32'hBE528484,
32'hBDE617FF,
32'h3F915FE5,
32'h3F18DE29,
32'hBF021A00,
32'hBE69CDA4,
32'hBEB9D308,
32'h3F0D349F,
32'h3F2BAFE1,
32'hBFC44D45,
32'hBF0C7F76,
32'hBF808331,
32'hBFB5F3C8,
32'hBE0AFE9E,
32'h3ED3C293,
32'hBF719877,
32'h3E97C5F2,
32'hBF17B2A8,
32'h3EA5ECEE,
32'hBD2AE533,
32'hBD89A91F,
32'hBF216301,
32'hBF7A059E,
32'h3F58BC4D,
32'h3F74576E,
32'h3EBD28E0,
32'hBF2F5921,
32'hBF8431DA,
32'hBD6D06FF,
32'hBEAFC825,
32'hBE1CB029,
32'h3DBB1E1C,
32'h3F180FF1,
32'h3EE478FA,
32'hBF5939CF,
32'h3DF335AE,
32'h3DD85326,
32'h3F2A6571,
32'h3E736340,
32'hBFFA1572,
32'hBF2CC308,
32'hBFA0CC0C,
32'hBFC244F2,
32'hBE47BF3A,
32'h3E67651C,
32'hBF73085F,
32'h3E9254E6,
32'h3E87457A,
32'h3F76E245,
32'hBD891489,
32'hBC113FEA,
32'hBD4179C9,
32'hBF2D83B9,
32'h3E918925,
32'h3EC43201,
32'hBD9C4252,
32'hBD23F815,
32'hBFCEAACD,
32'h3CEED740,
32'hBE909848,
32'h3E306D98,
32'h3EA3E619,
32'h3E426DD8,
32'hBEB2CFC4,
32'hBF14C5FE,
32'hBEBB8FE8,
32'h3D804995,
32'h3F6715DF,
32'h3E33AD61,
32'hBFD36023,
32'hBF2F2903,
32'hBFB9BE1E,
32'hBF72C9E3,
32'hBF1BA3EF,
32'hBEDF246A,
32'hBF78CE87,
32'hBEB86BCE,
32'hBE6C5292,
32'hBF904489,
32'hBE0BE2A2,
32'h3D3D5D59,
32'h2EC8BBFE,
32'hBEF54C09,
32'h3D7E6FD7,
32'hBEB59D93,
32'hBED76AFE,
32'hBEB44FF0,
32'hBF8CE435,
32'h3E1EC56E,
32'hBF86119C,
32'h3EC75D74,
32'h3EDC368C,
32'h3F7D47A5,
32'hBEB28A3B,
32'hBEFC9B2E,
32'hBF3197FC,
32'h3F296662,
32'h3F062E53,
32'hBE2D55A4,
32'hBFC05EA8,
32'hBEBD578B,
32'hBF96028D,
32'hBFD1DDAB,
32'hBF283DE7,
32'h3EF76FD1,
32'hBFF15FD3,
32'h3E33382E,
32'h3CB10B2A,
32'hBFE5785A,
32'h3D2421E3,
32'hBD4E714F,
32'hBE5B1E4C,
32'hBF54159A,
32'hBE01311C,
32'hBF0A5AD7,
32'hBFD2693B,
32'hBF3783EC,
32'hBFA43623,
32'hBF3CACFD,
32'hBF7D3253,
32'h3F174B1B,
32'h3E743DA1,
32'h3F5B4773,
32'hBEAAE2FE,
32'hBDACC42B,
32'hBE90A486,
32'h3F9B0035,
32'h3E6DFC68,
32'hBF18137B,
32'h3D091FBE,
32'hBDC1FE76,
32'hBEAA197F,
32'hBFF75B0D,
32'hBEE1BF95,
32'h3ECB2B59,
32'hBF98FFBB,
32'hBF27BBED,
32'hBE19E9DC,
32'hBF5F6043,
32'h3D22E4CD,
32'hBD412C48,
32'h3EFEE763,
32'hBF9B2835,
32'hBD75B6C1,
32'hBF655461,
32'hBFD30F7B,
32'hBED30F9B,
32'hBF9FF793,
32'hBE6810C2,
32'hBF924CA5,
32'h3F0A6905,
32'h3F73544D,
32'h3F90488E,
32'hBEE19ECF,
32'h3D3700BD,
32'hBF081774,
32'h3F453746,
32'hBE92CCC2,
32'hBF29ED3B,
32'h3E91FF99,
32'hBD39DA38,
32'hBF312C01,
32'hBEE27DC4,
32'hBEB3CA87,
32'h3E874464,
32'hBF00BCEF,
32'hBEAE1FF9,
32'h3F2E1A93,
32'h3DE65FB7,
32'h3C36DED2,
32'hBDF41EE7,
32'hBE490B9F,
32'hBF31428B,
32'hBDC323A7,
32'hBE7EAD0F,
32'hBFE53B81,
32'h5DE223C4,
32'hBFA59978,
32'h3DDE7E1B,
32'h3F0F06DD,
32'h3F13831E,
32'hBD82D8EE,
32'h3F21FD4B,
32'h3ED31C71,
32'h3D002BA1,
32'hBD8A619F,
32'h3EF60D47,
32'hBE868D6E,
32'hBE7CCDDE,
32'h3E36731D,
32'hBCF46E5D,
32'hBE58D89F,
32'h3E5E3FF4,
32'hBE8FF87F,
32'hBE2467B5,
32'h3E85875C,
32'h3D20CF30,
32'h3F17FE2A,
32'h3E03FA59,
32'hBD63BC63,
32'h3DC75926,
32'h3DAD88F0,
32'h3F8DD088,
32'h3F0F8B3A,
32'hBF6E7133,
32'h3F5E6351,
32'h3EC5F982,
32'hBF1F38FE,
32'h3E2245EC,
32'h3F37AE89,
32'hBE32DC6E,
32'h3E5E3321,
32'h3EA16D77,
32'h3F0F651B,
32'h3C76EB30,
32'hBCA5D81E,
32'h3EC8C3C5,
32'h3E5A03BD,
32'hBE3D0398,
32'h3DB6415E,
32'h5DD27249,
32'hBDA64EFB,
32'h3E3A0188,
32'hBE7BFEF9,
32'h3EAB90E5,
32'h3E6DE6DB,
32'h3E92A26A,
32'hBDC3704F,
32'h3EEBF840,
32'h3D113498,
32'hBC26367B,
32'h3E1BDA2A,
32'h3D398220,
32'h3D1CC697,
32'hBF273DF5,
32'hBD74081A,
32'h3F2E75AB,
32'hBDB2C389,
32'h3EAA2671,
32'h3E46385E,
32'hBD804F37,
32'h3DD9B1C7,
32'h3F1B28FD,
32'h3E053CFA,
32'h3C9946F1,
32'hBECFA68C,
32'h3EA19091,
32'hBDB3C310,
32'h3E96583A,
32'h3C6E132E,
32'h0ED345FB,
32'h3F7E2986,
32'h3D86895A,
32'hBDD41DA0,
32'hBF12547D,
32'h3F49D84A,
32'h3EEF1582,
32'h3F5211E2,
32'hBC5B696E,
32'hBCA5BAF0,
32'h3D3066C4,
32'h3E0A7C75,
32'h3EB8573F,
32'h3F79701F,
32'hBF922776,
32'h3E7EB643,
32'hBD9C8421,
32'hBE6300DA,
32'hBED18B79,
32'hBE3AA58B,
32'h3DC161B5,
32'hBD4A3525,
32'h3E175515,
32'h3EDC0D68,
32'h3D4576B4,
32'hBE7CCB84,
32'hBD9C8590,
32'h3F84B3B5,
32'hBE3CC699,
32'h3C120A16,
32'hBD7BB245,
32'hBA3BB39,
32'hBDAA09E5,
32'h5DF1B7C4,
32'hBE503D15,
32'h3F572612,
32'h5DCE411A,
32'h3F44E0CE,
32'hBD143E6B,
32'h3C8833DE,
32'hBD1002BC,
32'h3DCF314F,
32'h3ECC40CD,
32'h3C933036,
32'hBE8508BC,
32'hBD7523DB,
32'h3D4C68F7,
32'hBD5F85BB,
32'hBC785E10,
32'hBCA2E83C,
32'hBE9FBF7E,
32'hBD98E760,
32'hBE9F3FFE,
32'h3E833E91,
32'h1DF98D0F,
32'h3F106931,
32'hBD25EBD1,
32'h3F1A28DA,
32'hBC8888C9,
32'h3DAA758B,
32'hBCC05DCB,
32'hBCEC7826,
32'h0EDC0FC2,
32'h175053EA,
32'hBE8DAA3B,
32'h3F5EC4BE,
32'h3D29DAC7,
32'h3F444363,
32'h3C8B9F65,
32'hBDC2698F,
32'hBDB0DA3E,
32'hBE99591D,
32'h3F435775,
32'h3DF38F43,
32'h3D8537AE,
32'h3DDDBF7F,
32'h3C3180A5,
32'hBDBCAC75,
32'hBC967DBE,
32'h175AF4C1,
32'hBE2FEB17,
32'hBE5A416C,
32'hBF5E4A4A,
32'h3E3D1175,
32'hBDA282ED,
32'h3F4625F7,
32'hBDA1D70F,
32'h3F1F9AB0,
32'hBE893379,
32'hBDB4FBAF,
32'h3CDC8A6A,
32'h3D844526,
32'h3D98E837,
32'hBDB8089C,
32'hBCE3418A,
32'h3D7607B3,
32'h3DDD8AFC,
32'hBC9A08E9,
32'hBDE0AAF7,
32'h3DBA9B64,
32'hBCA892D4,
32'hBC086482,
32'h3CD51A0A,
32'hBCDC8510,
32'h3D215CB2,
32'h3D8C9CDD,
32'h3D4CF246,
32'h1DF1EEAF,
32'hBDC13550,
32'hBD00FD83,
32'hBD5C4F57,
32'h3C12F167,
32'h3CCA4DA5,
32'hBCBFA792,
32'h0EC4F7C5,
32'h5DF0442F,
32'h3DD5D65E,
32'h3CAC83B3,
32'h5DDC947E,
32'h3CCE5B7D,
32'h3D105C0F,
32'h5DDE36DE,
32'h3D4F8D5B,
32'h5DE0F447,
32'hBD2AA0A4,
32'h3C6DFE54,
32'hBCF7E19A,
32'hBD47EE8F,
32'hBD3D2383,
32'hBD3CE022,
32'h3D7C3A68,
32'h3DACC1FF,
32'h3C476566,
32'h3CF1CA10,
32'hBD3C2278,
32'h3DAF2C3A,
32'hBDA9AFEB,
32'h3C73F74F,
32'h1DCF1359,
32'h3DB73DD0,
32'h3D524A0C,
32'h3C16ED36,
32'h3D64364E,
32'h3DCD66EB,
32'h3DABD939,
32'hBC406728,
32'h3D84A8AA,
32'hBDCF0F75,
32'h3D690E81,
32'hBDCB6F6F,
32'h3D44DF7D,
32'h3D415E4F,
32'hBD4E6DE1,
32'h3CE5EC2D,
32'h0E5A460,
32'hBC07C03A,
32'h3CD60CF4,
32'h3DB380E2,
32'hBC6E7FFF,
32'h3D187320,
32'h3C7D03BB,
32'h3D06F676,
32'h3D0FECF2,
32'hBDD48BCA,
32'hBD80B170,
32'h3DA9FEFF,
32'h3D4F6A9A,
32'hBCD9F062,
32'hBC21BC16,
32'h3D348E67,
32'h3CC739C4,
32'h0ED060BC,
32'h3C203C09,
32'h3C8E58C8,
32'hBD0ABD24,
32'h1DF7E40E,
32'h3D8D5C84,
32'h3D32499B,
32'h3D22AC14,
32'h3C56394F,
32'h3D805A31,
32'h3D4AE6EB,
32'h3DDA8006,
32'h3D87B8D5,
32'hBC9CBB74,
32'h3CAA253D,
32'hBD1E0E86,
32'hBD0C2FB7,
32'h3D8BC46A,
32'h3D28FE96,
32'h3D988BE3,
32'h3D45E586,
32'h3D612E66,
32'hBC9F861D,
32'h3CF624CA,
32'h3D9094CC,
32'hBD8B41EF,
32'h07502932,
32'hBCCD8C07,
32'h3D1D8C56,
32'h3C1529D5,
32'h3D5FA168,
32'h3D61A280,
32'hBD7F3483,
32'hBC13C3A9,
32'h3D8D62E8,
32'hBCB15B8B,
32'hBD94A5C6,
32'h3D331128,
32'h3EE8BCED,
32'h0753F531,
32'h3DB98EFA,
32'h3C598394,
32'h1DC657F1,
32'h3D955FF7,
32'hBD1BA75A,
32'hBE2B2145,
32'h3D65CA6F,
32'h3F5467A6,
32'h3D8FD9AC,
32'hBC39B8D0,
32'h3D1208AB,
32'h3E056BDF,
32'h3D8F77C2,
32'h3F214826,
32'h3D88A1BC,
32'hBCB7D378,
32'h3DBD2A3B,
32'h1DDB68E0,
32'hBE2F0CEA,
32'hBEF73FCE,
32'hBF328225,
32'hBF5603D5,
32'hBE3CA2BE,
32'h3C9B28C5,
32'h3E113E77,
32'hBD134E8E,
32'h3D0CDD4F,
32'hBE9E9CE0,
32'h3F074058,
32'hBDC62FF4,
32'h3CB6AAA6,
32'h3DD6B7E6,
32'h3D9C4711,
32'h3CFF5509,
32'hBDEDE00E,
32'h3F136ECC,
32'h3DA7647D,
32'h3F33C5A9,
32'hBD6CE923,
32'hBCF3F725,
32'h3EA1220A,
32'h3E8EDD8D,
32'hBD17FEE0,
32'hBD6306AC,
32'hBD882C25,
32'hBECC616F,
32'hBE5508DD,
32'hBF2C15F8,
32'hBE52DCA0,
32'h3D117995,
32'hBF419788,
32'hBEBB29CD,
32'hBC2E9454,
32'h3D25E6A2,
32'h3F243DEB,
32'h3CB7688F,
32'h3D575767,
32'hBF76A587,
32'hBD6B1B15,
32'hBE206339,
32'h3E4E561E,
32'h3EC60633,
32'h3D5E1790,
32'h3E098D4E,
32'hBD85168E,
32'h3E85A0D7,
32'h075ECEF0,
32'hBD9E306D,
32'h3D5E93EC,
32'hBD92E128,
32'h3EDFBE0C,
32'h3C4000C2,
32'h3E055718,
32'hBF0907D8,
32'h3E121DF4,
32'hBE24A073,
32'hBEC5815F,
32'hBF2A9635,
32'h5DE8D7DA,
32'h3E000BA2,
32'h3D4953F7,
32'h3F3E6DF6,
32'h3E773D75,
32'h3DC84E84,
32'h3E84898C,
32'hBD29A8ED,
32'h3D70EA6E,
32'hBE5FBDAA,
32'h3CAE0599,
32'hBE27218B,
32'h3DC9CDC8,
32'hBEB5D301,
32'hBEA61138,
32'h3DD66CB3,
32'h3E6A3F96,
32'hBEA0544E,
32'hBDE67207,
32'h3E1A00CF,
32'h3D6CD667,
32'h3DBF9626,
32'h3E3DCE88,
32'h3C7F8E13,
32'h3DAE967A,
32'h3E9FEC11,
32'h3F07E869,
32'hBEE59835,
32'hBEEC5CE5,
32'h3E5AF521,
32'h3F43B1DA,
32'h3E6EE484,
32'hBE333003,
32'h3F12DD41,
32'hBEE6CBB7,
32'h3DDF2333,
32'h3E61AD2D,
32'h3E490D17,
32'h3D99BD60,
32'hBC0048C1,
32'h3CDD0F07,
32'hBD90B0A6,
32'h3ED49F97,
32'hBF5ABC1A,
32'hBDBC39E2,
32'h3D8B7F30,
32'h3F0DFD0D,
32'h3EC6DD64,
32'h3E4E3517,
32'h3ED64CAA,
32'h3D358B24,
32'hBC325F2B,
32'h3F0FF8F2,
32'h3F0423C3,
32'h3DB48CB3,
32'hBF39F20B,
32'h3F944458,
32'hBF3CA449,
32'hBF254EF5,
32'h3ED660D6,
32'h3E5181F9,
32'h3EA275B3,
32'hBE98710A,
32'h3F60A4FB,
32'h2EC13BFD,
32'hBC5B8C02,
32'hBE5F2F1A,
32'hBC5228F5,
32'h3F0A9527,
32'hBF0DBEC6,
32'h3F407D5D,
32'h3D250216,
32'h3F382158,
32'hBEC26582,
32'hBD9DD5E2,
32'h3E32682C,
32'h3F51C3BD,
32'h3F903A92,
32'h3EA6F09E,
32'hBEAAD073,
32'h3D9967BA,
32'hBCA54D0C,
32'h3E91BF2B,
32'h3FC2066D,
32'h3ED73914,
32'hBF03F59A,
32'h3E1CE812,
32'hBF824427,
32'hBF69D849,
32'hBEB68A5D,
32'h3E58B2A3,
32'h3EB5E807,
32'hBF1EFA20,
32'h3F03D5C6,
32'h3F02149C,
32'h3EA9F908,
32'h3EE0416C,
32'h3EA112EA,
32'h3E838D49,
32'hBF3BA517,
32'h3F1ABB0F,
32'hBDB5CEBC,
32'hBE4989A0,
32'hBF855B8D,
32'h3F37A8DE,
32'hBF1A5B09,
32'h3EF1C827,
32'h3F1A6011,
32'hBE31FC51,
32'hBE84FCF4,
32'hBDADD007,
32'hBD25DE5D,
32'h3D398996,
32'h3EA186FB,
32'h3DF1A7B1,
32'hBDB2634C,
32'hBD2D399D,
32'hBF4763BC,
32'hBFA33AFA,
32'hBEBAD1BB,
32'hBF1D716F,
32'h3F7D1813,
32'h3E8F19CD,
32'h3F9DD036,
32'h3DAEE229,
32'h3D809D88,
32'h3F42948C,
32'h3F25ABC0,
32'h3D96EA6A,
32'hBE9B5260,
32'h3F2777C1,
32'hBEC58220,
32'h3F05748D,
32'hBF57882A,
32'h3F476634,
32'hBFDB8882,
32'h3E94BB08,
32'h3F4C458C,
32'h3DC8A403,
32'h3F0D1075,
32'hBD424F75,
32'h3DAC2D41,
32'h3EC763EE,
32'h3F3BC983,
32'h3F058F68,
32'h3EA4333A,
32'h3F15C538,
32'hBF0301EE,
32'hBFB1E26C,
32'hBE8EDB79,
32'hBEEE2F49,
32'h3F4C537F,
32'hBF2516EF,
32'h3FBF537A,
32'h3CBC89E3,
32'hBD8CA825,
32'h3EB168A7,
32'hBE066ED1,
32'h3F5FD9F9,
32'hBD989B4A,
32'h3F349036,
32'hBF09F223,
32'h3F09C96F,
32'hBE90CCD3,
32'hBE9EFCC5,
32'hBFB7E8B7,
32'h3F3EB150,
32'h3F1F88A6,
32'hBEC780DC,
32'h3ED2FBCF,
32'h3DA41A72,
32'hBD322D6B,
32'h3E51C813,
32'h3EA700E6,
32'h3F1836E2,
32'h3E840734,
32'h3E36769B,
32'hBEAB7E28,
32'hBFEA40F1,
32'h3E70B396,
32'hBF145978,
32'h3F224D73,
32'hBF75E4AD,
32'h3FA221FC,
32'hBF239640,
32'hBF059B1F,
32'h3E642C6A,
32'hBEF52F7A,
32'h3F9881BD,
32'h3E9051D2,
32'h3E2C293C,
32'hBF3F81B6,
32'h3DB82683,
32'hBE0501FF,
32'h1DD05DC0,
32'hBFAD43C0,
32'h3F1C7EA4,
32'h3F235619,
32'hBE0FAE10,
32'hBEABAA3B,
32'h1DF1EE24,
32'h3CC07B63,
32'h3EA21D43,
32'h3EB0CC81,
32'h3F9957F3,
32'h3F41B50F,
32'h3E44722F,
32'hBE6039B1,
32'hBFF81FD9,
32'h3E1E1B42,
32'h3C94F525,
32'h3F1245AF,
32'hBF1DF0C9,
32'h3F976EFD,
32'hBEB6DAA7,
32'hBEB2D1C5,
32'h3F313AFD,
32'hBD80C659,
32'h3F514128,
32'h3EA27BDB,
32'hBE91906C,
32'hBE9F2B75,
32'hBF1AED97,
32'hBF233B32,
32'h3EB7964F,
32'h3DCC5AF0,
32'h3F86B8DA,
32'h3F9A6A1C,
32'hBF155075,
32'h3F62415B,
32'hBDBC6D6E,
32'h3CCA3EF1,
32'hBC5D2B29,
32'hBDE1A610,
32'h3D92A428,
32'h3EE58E23,
32'h3F229826,
32'hBD71250F,
32'hBF9581F2,
32'h3D936A05,
32'hBF006CEA,
32'h3E9C86CD,
32'hBF7CED24,
32'h3F5EF85F,
32'hBF0FC273,
32'hBEC58459,
32'h3F52844F,
32'h3E1568F8,
32'h3DF3A4BE,
32'hBE8A4CD8,
32'hBF5A7D44,
32'hBF026B4B,
32'hBEB1239D,
32'hBF38C6B6,
32'h3E13E927,
32'h3F388B92,
32'h3EBB1E7E,
32'h3F635D1A,
32'hBF70959D,
32'h3F1764F9,
32'h3C737AAB,
32'h3D22C305,
32'h3F27D9A0,
32'h3E82503E,
32'h3ED4E9E4,
32'h3E80A5A0,
32'h3F0B4C9A,
32'h3DD352CB,
32'hC040F51E,
32'h3C23DBE4,
32'hBF6FFFD7,
32'h3E161F53,
32'hBEE5B7B9,
32'h3F2E47E8,
32'hBED2BDA6,
32'hBF0211CD,
32'h3E63DA5B,
32'hBEB180FD,
32'h3ED9E973,
32'hBEE8FC20,
32'hBFF4716D,
32'hBF2B6D63,
32'hBF051C1A,
32'h3E1EAA34,
32'h3EE4D75F,
32'h3CFDD95E,
32'h3E85B70A,
32'h3F6C1FA5,
32'hBEE7DD41,
32'h3D1D8825,
32'h3C7E8CE6,
32'hBD149B1D,
32'h3DF9CD86,
32'hBE64E0DB,
32'hBE5B00E3,
32'h3EB5B376,
32'h3EE84E03,
32'hBE9519E0,
32'hBF73633A,
32'hBD8C87BF,
32'h3C9BB808,
32'h3E8001D5,
32'hBD2813D8,
32'h3F546CF2,
32'hBE1280B0,
32'h3EFEFD5F,
32'hBD4EB6D2,
32'hBDA697B4,
32'h3F458B66,
32'hBE3FE6D3,
32'hBF925AA8,
32'h3EEAE827,
32'hBE342EC6,
32'hBE723AD0,
32'h3EF458ED,
32'h3ECA986E,
32'hBEEE2BB8,
32'h3F432DBA,
32'hBE9B45EA,
32'h3F4A05C1,
32'hBD957605,
32'hBCE8A816,
32'h0EDE11AE,
32'hBE031978,
32'hBEB82556,
32'h3ED76A5F,
32'h3E9F7673,
32'hBF269C41,
32'hBFB56316,
32'hBD78F3F6,
32'hBF93250C,
32'h3D9208ED,
32'hBE41DC28,
32'h3F3310D0,
32'hBE1C5A44,
32'h3EB0FD00,
32'h3DAC777E,
32'h3E30AF8A,
32'h3F13840B,
32'hBE80316D,
32'hBEAD0EA5,
32'h3E81AABD,
32'hBF25777D,
32'h3EB6868A,
32'h3EFBDC0A,
32'h3E0C151A,
32'hBF1804BD,
32'h3F51553B,
32'h3EA44970,
32'h3F157DC7,
32'h3D8363EC,
32'h3D721870,
32'h3E40E112,
32'hBDB0F4F1,
32'h2EC4DE19,
32'h3E773A7A,
32'h3E24FB74,
32'hBF09205A,
32'hBF288E7A,
32'h0ED24E76,
32'hBFBCAA76,
32'h3EA921C7,
32'h3DDF6DE1,
32'h3F2ADFAA,
32'h3DA5447C,
32'hBE0AF679,
32'hBE96C10B,
32'h3F13437C,
32'h3F1963FA,
32'hBE2F8223,
32'h3E064009,
32'hBCBEEB81,
32'hBF2EB614,
32'hBEE1E3F1,
32'h3DC0E6BE,
32'h3EBAAAEF,
32'h3ED2B21B,
32'h3E569A0E,
32'h3E93FFE6,
32'h3E678F08,
32'hBDA45BDC,
32'h3D25D135,
32'h3E5D6C72,
32'h3C6B42A4,
32'h3E94E7B8,
32'h3ECA5C8E,
32'h3DCA8A8C,
32'hBEC45AEF,
32'hBDB5371F,
32'hBD9DBBC4,
32'hBECC6EDF,
32'h3DD81674,
32'hBD9DC42E,
32'h3F2501BA,
32'h3E8C7F72,
32'hBE9FE705,
32'hBE1548D2,
32'h3EE0AE49,
32'h3F7218E0,
32'hBE31E12B,
32'h3EB4C418,
32'hBDF4F27F,
32'hBF90FA9C,
32'hBF244516,
32'h3D8908B5,
32'h3F3D5893,
32'h1DE29596,
32'h3EFE481F,
32'hBE0765FC,
32'h3E3676C6,
32'h3DB07A04,
32'h5DF7010E,
32'hBDC2BF9B,
32'hBCBFF91B,
32'h3F075813,
32'h3DA5A85D,
32'hBD00376F,
32'hBEC6AFFB,
32'hBEEE0F92,
32'hBDE6B7DA,
32'hBF3EF0FA,
32'h3E8EDE99,
32'hBE361058,
32'h3F50ABC8,
32'h3EF55C5D,
32'hBE99ED9E,
32'h3D70ACA5,
32'h3F2CDD6D,
32'h3EDE52F6,
32'hBE600B99,
32'h3E78BF5A,
32'hBDAE5F7B,
32'hBECF1EC7,
32'hBF33F4FE,
32'h3EE194AD,
32'h3DD09783,
32'hBE1CDF09,
32'h3E50D6E5,
32'hBDE1BF76,
32'hBEE172EF,
32'hBD934FCE,
32'h3C96B23F,
32'hBE0C4D3A,
32'hBEA4A9B4,
32'h3F3D796F,
32'hBD431743,
32'h3ED0B51E,
32'h3DF8FDA6,
32'h3E925488,
32'h3F2F29AA,
32'hBEEF381F,
32'h3D874091,
32'h3E105F54,
32'h3F551534,
32'hBED95056,
32'hBE1F8993,
32'hBEE323F6,
32'h3EFCE9D0,
32'hBCC5A178,
32'h5DFDEB79,
32'h3ECA40B9,
32'hBE4B81E6,
32'hBF94865C,
32'hBE5E6398,
32'h3EAC2DA1,
32'h1DCA203C,
32'h3EABB093,
32'h3F8E91DB,
32'hBEECFE01,
32'hBF1400AB,
32'hBCB05CAE,
32'h3DB17FF7,
32'hBEC78F79,
32'hBEFF7634,
32'h3E36BAC0,
32'hBDFF627A,
32'hBEAAB784,
32'hBDB42FDA,
32'h3ED07A6B,
32'h3E6A1222,
32'hBEE5EBFE,
32'h3EC5198E,
32'h3C5EF218,
32'h3D3B9725,
32'hBEBF90D0,
32'h1DC67840,
32'h3E6A281D,
32'h3F53A344,
32'h3EC4845F,
32'hBF2C25CE,
32'h3D9C81AB,
32'hBE3065A3,
32'hBF2B68E5,
32'hBE631E75,
32'h3F574D70,
32'h3E94456A,
32'hBF95A9A1,
32'h3E8866FE,
32'h3D7F231C,
32'hBF469294,
32'hBD10042F,
32'h3CCF150F,
32'h075349D0,
32'hBF2B001F,
32'h3EF4DED1,
32'h175CF8A3,
32'hBEF53719,
32'h3EE7197F,
32'hBF02C650,
32'h3ECF2EE6,
32'h3F325FC7,
32'h3F232EE1,
32'h3E03D8DD,
32'h3EF7F781,
32'h3D19B84C,
32'hBD519392,
32'h3D31BA0F,
32'h3EBDDC91,
32'h3E436ED7,
32'hBF07453C,
32'h3ECABFEB,
32'h3D0760FD,
32'h3D7A8B10,
32'hBF26FE94,
32'h3F423CED,
32'h3DA265C7,
32'hBFA5A922,
32'hBE8D8B7E,
32'hBDACE00F,
32'h3F8FDCEA,
32'hBDD87271,
32'hBC26FE38,
32'hBE888F61,
32'h3F2CB247,
32'hBDBA3CC8,
32'h3CF44069,
32'h3F3046D3,
32'h3EEB928C,
32'hBFB3BFB9,
32'h3EFE744B,
32'hBD1845F2,
32'h3D0EA8C6,
32'h3EC02921,
32'h3EB0CDB9,
32'h3EB558FB,
32'h3E71894E,
32'h3EC5C474,
32'h3C5D7CD7,
32'h3D8D9E3B,
32'hBD85D8D4,
32'h3EACC971,
32'h3EE657F3,
32'h3F72CC75,
32'hBE32ACF2,
32'h3F033289,
32'hBE02EE65,
32'hBFCFBB77,
32'h3F28BEBE,
32'h3DEFE45E,
32'h3C7FA154,
32'h3DD2417E,
32'hBD885B69,
32'hBEB3D0E5,
32'hBF08379D,
32'hBEA78EE2,
32'h3E97645D,
32'h3EB9203B,
32'h3E5A1854,
32'hBCF42F8F,
32'hBEBBF489,
32'hBE9592E7,
32'hBD5EF0D0,
32'hBF96BA13,
32'h3F75FBF6,
32'hBF133EDD,
32'h3C51D19D,
32'h3D3793ED,
32'h3D031E29,
32'h3D4DFDE2,
32'h3E6720F3,
32'hBEB4E1CB,
32'h3EBB2757,
32'hBD1043E6,
32'hBE066B40,
32'h3E5CDA46,
32'h3ECA090D,
32'hBF079CA0,
32'h3EA39974,
32'h3ED8E517,
32'hBD990F91,
32'hBCB12949,
32'hBC0871A3,
32'hBF0929C4,
32'hBDE65E45,
32'hBF1A6EBB,
32'h3E6E5581,
32'hBE58D93D,
32'h3EDC2C17,
32'h3D5C7769,
32'h3DCC43B5,
32'hBEA26B1E,
32'h3F21B5A2,
32'hBF685DBD,
32'h3D30717A,
32'hBE83FC3D,
32'h3D8DF95A,
32'h3E873B8D,
32'hBD29BEA0,
32'h3E8103E6,
32'hBF00D91B,
32'hBEAC8220,
32'h3D8BB51A,
32'h5DE9CE33,
32'h3EBBCEC0,
32'h3D1947EF,
32'hBEBC9CD7,
32'h3E6BC499,
32'h3EBF9FD0,
32'h3F227935,
32'hBDC28F9A,
32'hBD938A2F,
32'h3D49E406,
32'hBD8B04F7,
32'h3F1BAAD7,
32'h3DE34FB4,
32'h3E108CD8,
32'hBDDB7751,
32'h3E2165D8,
32'h3DCF28C2,
32'h1CF4EAA,
32'h3DB4F453,
32'hBEF13218,
32'hBEB2837E,
32'hBE358F7A,
32'h3DB5A56A,
32'h3C6141DA,
32'h3D9D914A,
32'hBEFDB28C,
32'h3EF9856A,
32'h3E9181A4,
32'hBE30023A,
32'hBD01BBBE,
32'h3DC7B6B9,
32'hBCF1BC24,
32'h3CF7C2E2,
32'hBD788C5E,
32'hBD69DC44,
32'hBDD7067E,
32'h3D0FB3D0,
32'hBD984C27,
32'hBD7EBDF6,
32'hBC18062F,
32'h3E67D442,
32'hBDCE07DB,
32'hBCAACAB4,
32'hBE84EC8E,
32'h3D050351,
32'hBC30F3B4,
32'hBC0813C5,
32'h3D286BEF,
32'hBD983F0C,
32'h3E6B68B8,
32'h3D239362,
32'h3EDD123F,
32'hBDBB50DD,
32'h3D1242D1,
32'hBE92D58C,
32'h3C6346A0,
32'hBDCCABDC,
32'h3E93C64A,
32'h3D6B5811,
32'hBD57AD57,
32'h3C588090,
32'h3D2C474F,
32'hBD4E3B2B,
32'hBC169125,
32'hBCE68F00,
32'hBCA74B62,
32'hBD1B5E2B,
32'hBD7D9DDA,
32'hBC947D31,
32'h075C438E,
32'hBCE17117,
32'hBDC13B26,
32'h3C1B705D,
32'h1DE23F88,
32'hBC963135,
32'h3C2050B3,
32'h3CDB97E3,
32'h3DC6A4FA,
32'hBD0E9D33,
32'h3D264AB2,
32'h3D52A015,
32'hBCA47D2A,
32'h3D503548,
32'h1DF51BE9,
32'h2ECAFE67,
32'h3CE7237C,
32'hBC842A67,
32'hBCEF426D,
32'hBDCFC25D,
32'hBC73FD53,
32'hBD8CEEEF,
32'h3CCC17E0,
32'hBD32D488,
32'h3D7890F6,
32'h5DE98C82,
32'h3D8C501F,
32'h3C613BA3,
32'hBC626BFA,
32'h3D9C7C9D,
32'h3CC24F90,
32'h3D5D148B,
32'hBDD74259,
32'h3D246FE4,
32'hBCA13D5B,
32'hBD118F27,
32'hBD04FBE0,
32'hBCACD15D,
32'hBC31FA09,
32'h3D81EC8C,
32'h3D74BC88,
32'hBCFC9ED3,
32'h1DD11871,
32'h3C0ED4A9,
32'h3D0CB3C7,
32'h5DE1F867,
32'h3DCA1002,
32'hBD9B1F6F,
32'h3D28A24A,
32'h3D003252,
32'h2EDC6BAB,
32'h1DC445C5,
32'hBD15D13C,
32'hBD4BEF79,
32'h3D41875F,
32'hBEC3BF1A,
32'hBD3A0F70,
32'h3D7177A0,
32'hBD04325A,
32'h3D199BEA,
32'hBD814C09,
32'h1DF8F5C4,
32'hBD89A0AB,
32'hBCB3BCA6,
32'hBEA798D9,
32'hBDB751D6,
32'h3D7BAA27,
32'h5DEB585F,
32'h175B8DD9,
32'h3C108F6A,
32'hBE2A4EFF,
32'h3CF8E9B1,
32'h3EE44116,
32'hBF0ECEB5,
32'h3D8A4C3E,
32'hBF045F3C,
32'hBCB9B459,
32'hBE2905FC,
32'h3E01DE07,
32'h3ED8817F,
32'h3DC63FC2,
32'h3DF649B4,
32'h3D189618,
32'h3D3469F4,
32'h3D8D2D62,
32'h3E50288D,
32'h3E889CB2,
32'h3CDDA96A,
32'h3F385336,
32'h3C6C7DD3,
32'hBA3E976,
32'hBE0D02E1,
32'h3E2E05AD,
32'hBD33AC8B,
32'h3F51D7D8,
32'hBCCE9AA7,
32'hBC6FA00F,
32'h3C7B2B48,
32'hBC177320,
32'hBE663A05,
32'hBF33CE3D,
32'hBF2D6F0D,
32'hBF828DCA,
32'h3D495FC8,
32'h3D4FAF2E,
32'h3E4EABDA,
32'hBD672299,
32'h3DA5B5A2,
32'hBEAF2001,
32'h3EC7E0C8,
32'hBCE57BDA,
32'hBEAEFA94,
32'h3E59CD6D,
32'hBE029652,
32'h3CD499ED,
32'hBE6BF4BB,
32'h3F48A42B,
32'hBD9E12EF,
32'h3F38123D,
32'hBD6FC929,
32'hBD2B7886,
32'h3C88AD4D,
32'hBEAC2754,
32'h3E12E28D,
32'h3F26A534,
32'hBD87D3DF,
32'hBF09B162,
32'h3E83DFFB,
32'hBE8F05A3,
32'hBDAB5B01,
32'h3F209572,
32'hBF293092,
32'h075B0089,
32'hBF04566E,
32'h3E9FD5F1,
32'h3E086B05,
32'h3E9FCD0C,
32'h3E199E1B,
32'hBF80F0B1,
32'hBE88A266,
32'hBEAD0C38,
32'h3E386B37,
32'h3EC6DCE2,
32'h3F10BBC2,
32'hBEBA4E8D,
32'h3F499665,
32'h3E3D04EA,
32'h3E9FADB3,
32'hBCDEA8BC,
32'h1DD9E408,
32'hBC9325EB,
32'hBF9FA39D,
32'h3E4895DC,
32'h3F17ECFB,
32'hBE8F9C42,
32'h3EC77164,
32'hBE3277A7,
32'hBF0FB15F,
32'h3E1F23FA,
32'h3E1D5912,
32'h3EDB6B56,
32'h3C88FE76,
32'h3F1B488E,
32'hBDB02C54,
32'h3E127620,
32'h3F22EC14,
32'h3F39EACA,
32'h3E94FB54,
32'h3DF40726,
32'hBE836096,
32'h3DEC5406,
32'h3DC8366D,
32'hBF28D19D,
32'h3F0FB496,
32'hBF19D854,
32'h3FA8BC3E,
32'h3E9EB816,
32'h3DFD2D0C,
32'h3F32C845,
32'hBC515CC7,
32'h3D1010DE,
32'hBF8903D6,
32'hBEFB40BC,
32'h3F33CDB0,
32'h3E1C31E0,
32'h3F160E17,
32'h3F3D7A32,
32'hBCB3C3B4,
32'h3F434AB0,
32'h3F135CBC,
32'hBE7C7985,
32'hBE559F57,
32'hBF409670,
32'h3F62B597,
32'h3F1D0CC3,
32'h3EFE0BF5,
32'h3F564793,
32'h3DCC34C1,
32'hBE8A89F2,
32'hBE411094,
32'h3EC69F43,
32'h3EB884E8,
32'hBF336CA4,
32'h3F03B8BE,
32'hBF88C270,
32'h3F359C51,
32'h3EA587AD,
32'h3F1F62DF,
32'hBE3647FC,
32'h1DC6F1C8,
32'hBC0F6A61,
32'h3D71825E,
32'h3E611198,
32'h3EB04012,
32'hBF09B262,
32'hBC995252,
32'h3E68E7BE,
32'h3D80EE9A,
32'h3E326E05,
32'h3E85801C,
32'h3E744ABE,
32'hBEE499E8,
32'hBE888C98,
32'h3F0C4876,
32'h3F3DECD7,
32'h3D623B7C,
32'h3F34EAFA,
32'h3CADEC3F,
32'hBF88FB0F,
32'h3F3A6A9E,
32'hBF93D6D6,
32'h3F20618E,
32'hBEE8663C,
32'h3F237A26,
32'hBFAB021A,
32'h3CAE4718,
32'hBE0BF939,
32'h3E684E4C,
32'h3F1804A8,
32'h3D09D078,
32'hBD54C4A3,
32'h3DBC4587,
32'h3F06A258,
32'h3EA3B197,
32'hBCA7B001,
32'h3F3BEF26,
32'h3F56A1A1,
32'hBDD319BF,
32'h3E393D6A,
32'h3F0FA5D5,
32'h3F003ADB,
32'hBFB8722F,
32'hBEA87179,
32'h3F135882,
32'hBF075775,
32'hBCC5C547,
32'h3EB4493A,
32'hBE5EF861,
32'hBF25266C,
32'h3EEDC9CB,
32'h3E81EC96,
32'h3EE5B650,
32'hBE32C0FF,
32'h3F7126AE,
32'hBF6107CF,
32'h3F694A0F,
32'h3D709145,
32'h3F239150,
32'hBE269214,
32'hBD86F83C,
32'h0754CAF0,
32'h3EA8DAAE,
32'h3DD59A99,
32'hBEEE76E1,
32'h3EA450FD,
32'h3E45D650,
32'hBE8A2D70,
32'hBEEA50B2,
32'h3D903FA8,
32'hBE65F054,
32'h3EA5E60E,
32'hBEB1721F,
32'h3ED73D74,
32'h3EB1EAF4,
32'hBE2F0D6B,
32'h3D831771,
32'h3EB446EF,
32'h3E617B88,
32'hBF12E51E,
32'h3EAF9CE2,
32'hBDAB9276,
32'h3E258F8F,
32'hBEBC2D53,
32'h3E899487,
32'hBC58A35E,
32'h3E789FE8,
32'h3E150232,
32'hBE899F8A,
32'hBF28A645,
32'h3D34DF62,
32'h3D2ED010,
32'h3EB1CEDA,
32'h3ECC08B8,
32'hBE24BB8F,
32'h3EC270EE,
32'h3E0F3C2F,
32'hBE92E510,
32'hBF981C72,
32'hBC605A4D,
32'hBEABF692,
32'h3EBC4201,
32'h3CA9570F,
32'h3F020877,
32'h3ECC6123,
32'hBF40512E,
32'h3D5BA9E4,
32'h3E63BA3C,
32'h3EDFDEB1,
32'hBE01E961,
32'hBEFA4A0D,
32'hBF091085,
32'hBE86F288,
32'hBE8899A6,
32'hBF7A50D5,
32'h3ED28349,
32'h3F0044E0,
32'h3EBB9B1E,
32'hBE2DDAAB,
32'h3E4A8239,
32'hBD94ABC0,
32'h3D15972A,
32'h3F03DF5C,
32'h3EE98217,
32'hBE8EF961,
32'h3DF60FAC,
32'h3D12755C,
32'hBD980080,
32'hBF3A374E,
32'h3DE24BC8,
32'hBF189AC7,
32'h3DC93647,
32'hBF0EDD3D,
32'h3D9431C4,
32'h3E3D35BF,
32'hBF1DC298,
32'h3E881BC2,
32'hBE295EBE,
32'h3E68C7EF,
32'hBE82FD28,
32'hBECDC9FC,
32'hBEBADA00,
32'hBECEEC8F,
32'h3DEE7904,
32'hBF606186,
32'h3ECD398A,
32'h3EF695E3,
32'h3E3BEAEB,
32'h3EB6F5E5,
32'h3EB0BDEF,
32'h0ED6982E,
32'h3D893E18,
32'h3EA87550,
32'h3E9D8EAD,
32'hBE7DEF7C,
32'h3E1CE810,
32'h3F0D3E78,
32'h3E69C9F0,
32'hBE8295AE,
32'h3E86A56D,
32'hBF125C80,
32'h3E182C81,
32'hBF44AC53,
32'hBE13444E,
32'h3EB9468B,
32'h3E1CC641,
32'h3EBA5F4A,
32'hBEAF9143,
32'h3EDE2A93,
32'hBF1C3C2F,
32'hBEA7BDFB,
32'hBE701C3F,
32'hBDA72345,
32'hBE2FB6E7,
32'hBF3FD0A3,
32'hBE150AA3,
32'h3EDC5CF7,
32'h3E36EBCE,
32'hBE3DE130,
32'h3CF8C205,
32'h3D3E2DA8,
32'hBCE7B1B7,
32'h3C20387B,
32'h3F20B09B,
32'hBE58D355,
32'h3E94A23D,
32'h3F07AAF7,
32'h3E2DC488,
32'hBCBD6888,
32'h3EE2165C,
32'hBF093DA0,
32'h3E33EADA,
32'hBEEA9BC2,
32'h2ED6B30D,
32'h3CE4EBD2,
32'hBE418EB8,
32'h3E6F8823,
32'hBEFFCBC9,
32'h3E1A6A86,
32'hBF0C5CFE,
32'hBF79B7E9,
32'hBE5BA880,
32'h3EC72AA3,
32'h3E143F91,
32'hBE8C87DF,
32'hBE0628C4,
32'h3E214690,
32'h3E49B9F8,
32'hBF78B1F0,
32'h3DE60492,
32'hBCA8FC00,
32'hBD111D51,
32'h3D939405,
32'h3E42A9E6,
32'hBE99844A,
32'h3E685C2E,
32'hBD2132D2,
32'h3E216CD2,
32'hBF145D15,
32'hBD470D7D,
32'h3D2FF62A,
32'hBD3CD1B1,
32'hBEFCBD24,
32'hBDD12051,
32'hBE9C5C89,
32'hBEEC661E,
32'h3DF46676,
32'hBE4A8FE6,
32'h3DEBD9B5,
32'hBEBC542C,
32'h3D5EE7FC,
32'hBEA5ACF8,
32'h3E324A4D,
32'h1DC96BE0,
32'h3D35A2E4,
32'h3D833E4F,
32'hBC0E485F,
32'h3E41349D,
32'hBF7AEFFB,
32'h3C3BAB34,
32'h3D5B7F6F,
32'h3DB9F7F3,
32'h3E43C340,
32'h3E38AC9B,
32'hBDF0768E,
32'h3E19BEE9,
32'h3DAC4D3C,
32'hBF357149,
32'hBFB8D8E0,
32'h3E9E9140,
32'h2ED8B274,
32'h3DA64605,
32'hBE87289B,
32'hBE0B940B,
32'hBE484936,
32'h3EE87039,
32'h3E9A1F86,
32'hBE53A1F5,
32'h3E6AAAA2,
32'hBED69381,
32'h3F5D6539,
32'hBF1004F3,
32'hBD00B8F5,
32'h3D04152D,
32'hBEFD9A5B,
32'h3DD55DE9,
32'h3DA7B2BA,
32'h3E497450,
32'hBF22F8AC,
32'h3E114C6A,
32'hBE1B44CE,
32'h3C85F6E1,
32'hBDE6E79C,
32'h1DC30C82,
32'h3DED9C38,
32'h3E06AEF2,
32'hBEA22DC4,
32'hBF7E38B8,
32'hBF8CB9E4,
32'hBEB2EBE2,
32'hBF1CEA35,
32'h3E4DEB74,
32'hBE089F1B,
32'hBE3321FD,
32'h3D92C248,
32'hBE355F14,
32'h3E2D5FC4,
32'hBE790E2B,
32'h3E9ADCB8,
32'hBE36A975,
32'h3E88D35F,
32'hBD073A33,
32'hBE4898AE,
32'h3E6E0467,
32'hBF3CC0F6,
32'h3C0CE3BC,
32'h3E105CB7,
32'hBC1AF71A,
32'h3D8C238C,
32'hBE23EC4E,
32'h3C9C7068,
32'hBD8EBF3B,
32'hBEA9473E,
32'hBD6542D3,
32'h3E050385,
32'h3E210ACA,
32'h3E90AAF9,
32'h3CF928BE,
32'h3C29EF33,
32'hBECAD1C2,
32'hBCEBF2DE,
32'h3E7A9D4B,
32'hBE20CC36,
32'hBDD0BBBF,
32'hBE004436,
32'hBEAF9777,
32'h3D9E090F,
32'hBDD9879D,
32'h3EDBB6E3,
32'h3E38EDCA,
32'h3E1FE441,
32'hBE4C9832,
32'hBE7F2B02,
32'hBD8EAC25,
32'hBF4F8479,
32'hBD628878,
32'h3E242770,
32'hBE849B5D,
32'h3E8F9195,
32'h3E52E7F0,
32'hBDA446EA,
32'h1DE970B8,
32'hBE74B298,
32'h3E870441,
32'hBE0C7604,
32'h3DC59A92,
32'hBD0009EA,
32'hBEFAE1E3,
32'hBEEB4B28,
32'hBDA97CD5,
32'h3CBF889E,
32'h3E89D4B3,
32'h3E4DBB41,
32'h3E0F47D4,
32'h3D279B63,
32'h3D80EB42,
32'h3E127F42,
32'h3E2FC8F1,
32'h3F08D80D,
32'hBE8648DF,
32'h3E5AE81B,
32'hBEB38B01,
32'hBDFA207E,
32'h3EEBA15F,
32'hBE75B0B9,
32'h3EC8436F,
32'h3DD1701C,
32'hBD61C901,
32'hBDBAA92B,
32'h3DD84172,
32'hBCC49524,
32'hBDD0D8B5,
32'h3C54B93B,
32'h3E94DB20,
32'h3D876FD4,
32'hBE9AF8CD,
32'hBE0C20F3,
32'hBE660FF8,
32'hBEBC6071,
32'hBEF959AE,
32'hBECC7778,
32'h2ED59E0A,
32'hBED881F8,
32'hBD413AD0,
32'h3D9162DF,
32'hBF8356FC,
32'h0EDEF38D,
32'hBDE72737,
32'h3E9559D7,
32'h5DFE10C1,
32'h3F0CF4A2,
32'h3EB3A1C3,
32'hBEA36C3C,
32'h3D70E93E,
32'h3EB7D9AC,
32'h3D294450,
32'hBE3C73C5,
32'hBE286FDE,
32'hBE30492E,
32'hBF027BAD,
32'hBC138101,
32'h3C941642,
32'hBED3C67D,
32'h3E361D9E,
32'hBDEEB77A,
32'h3CC1A858,
32'h3EE2B92A,
32'hBDBA89E7,
32'h3EEF59CA,
32'hBD48F6E2,
32'h3ED9C29C,
32'hBE9354F4,
32'h3E50CA3E,
32'hBE7F25A6,
32'hBD992A61,
32'hBE5256CA,
32'h3CF4B7F6,
32'hBE8D8BC3,
32'h3D5E5F84,
32'h3D92D1EB,
32'h3F33C96B,
32'h3D31FFD7,
32'h3E90C863,
32'hBE4D701C,
32'h3F2AAAC1,
32'hBE6E06F9,
32'hBEC4E92B,
32'hBC9818DA,
32'hBE981F62,
32'hBF4014EC,
32'h3DAC2A68,
32'hBCCE57DC,
32'hBED96570,
32'hBD78B012,
32'h3DCC0A39,
32'h3E0E7682,
32'h3DE10A0E,
32'hBDA32059,
32'h3E8DF6C0,
32'h3E635E88,
32'h3E2F2AC9,
32'hBC1C26F5,
32'h3EDF888B,
32'hBD3EB8B3,
32'h3D0B2BA4,
32'hBEDB5988,
32'h3E2654AB,
32'hBE14C737,
32'h3D08F1E1,
32'h3E1E5CEF,
32'hBDC9AD68,
32'h3DEEFF84,
32'hBE441E4B,
32'h3D9A5411,
32'h3F863B4C,
32'h3E5FEE2B,
32'hBF014428,
32'h3D3E9538,
32'hBEE74AC0,
32'hBF296707,
32'hBD96B34B,
32'hBD1CF16E,
32'h5DC48E94,
32'hBEABEB58,
32'hBE49BD41,
32'h3C3E3E56,
32'hBF293750,
32'h3F19FAD4,
32'h3E75721C,
32'h3EC78412,
32'h3EA3998E,
32'h3F080B3E,
32'hBDEDD3E0,
32'h3E28ED83,
32'hBECEF980,
32'hBEBCED8A,
32'h3EC7949B,
32'h3DA8372A,
32'hBD27468A,
32'h3EF36805,
32'h3EE4921D,
32'hBE2FFEC1,
32'hBE2543EA,
32'h3E1B53F5,
32'h3F9E3958,
32'h3EC2D538,
32'hBECE388B,
32'hBDCC45AA,
32'hBEFE4574,
32'hBEBF2CF9,
32'hBD15ECB0,
32'h3CACC571,
32'hBD771582,
32'h3EAB76EC,
32'h3E8C90D3,
32'hBE3F261D,
32'hBE2F11F7,
32'h3F60DE3D,
32'hBC707B42,
32'h3F52DC3B,
32'hBED1F335,
32'h3DB33F0B,
32'h3DE97ADD,
32'h3E5A7250,
32'h3F039F39,
32'hBEED1A79,
32'h3EFA94A0,
32'h3E19FA00,
32'hBEBA4C22,
32'h3E78B8CB,
32'h3CB81C2B,
32'h3E35A403,
32'h3F161D87,
32'hBE2D6F07,
32'h3F5C9F2C,
32'h3F0F5799,
32'hBEC2AFD2,
32'hBE83E17A,
32'hBED8390E,
32'hBF12D9E6,
32'h0ECD3974,
32'h3CCF6256,
32'h3D88B938,
32'hBF346714,
32'hBF0ACCA3,
32'hBE710AD6,
32'hBEA43102,
32'hBE4AD751,
32'h3E7FF6BD,
32'h3F2443DE,
32'h3F266082,
32'h3EC1A9A2,
32'hBE0635CD,
32'h3EB24257,
32'hBF6CDCAE,
32'h3D87408F,
32'h3F2109D5,
32'h3EB933CD,
32'hBE867027,
32'h3E12A87B,
32'hBF15D23C,
32'h3EE10750,
32'hBEB9C4C7,
32'hBE53F70C,
32'hBD11175F,
32'h3EA274C0,
32'hBEAA933F,
32'hBD57341A,
32'hBED1F0F6,
32'hBE3596B6,
32'hBD0A0CB8,
32'h3C22B9B0,
32'hBE373205,
32'hBFABD716,
32'hBFBDA1A8,
32'hBF31AC9B,
32'hBF2A8F48,
32'hBE8C40AD,
32'hBE99B3E9,
32'h3EADD15E,
32'h3ED5ACBA,
32'h3F753898,
32'hBFC18F19,
32'h3EAB7324,
32'hBEDFFA30,
32'hBD46CF76,
32'h3F7285F6,
32'h3EE2702F,
32'hBEFE3A35,
32'hBE9F1A77,
32'hBF65B36D,
32'h3F083024,
32'hBF469FAD,
32'hBF04371F,
32'h3F905311,
32'h3ED62D1A,
32'h3EEA1974,
32'hBEBBE44F,
32'h3F4515F0,
32'h5DEE7EEF,
32'hBCB1DE19,
32'hBDD5FECA,
32'h3E394E97,
32'h3E52F71B,
32'hBF81E3B7,
32'hBED44FA5,
32'hBF93A0C9,
32'h3F09FFE0,
32'h3F812003,
32'h3F8D284A,
32'h3E3E0807,
32'h3EF49BB6,
32'hBED91F88,
32'hBED3C532,
32'hBD417F02,
32'hBD565E8A,
32'h3F2CED5B,
32'h3F0CDF26,
32'h3EA4178F,
32'hBF7A0719,
32'hBE7523FD,
32'h3C657365,
32'hBE3F33E5,
32'hBE9FFE78,
32'h3F077BB7,
32'h3F36BA93,
32'h2ECDB585,
32'hBEDE004A,
32'hBCDF69EF,
32'h3D2DDEDA,
32'h3D101576,
32'hBD2DB8CE,
32'h3EA068BE,
32'hBD82A2F2,
32'hBE019404,
32'hBCFDB00F,
32'hBF057AA6,
32'h3E50D86F,
32'h3D31008F,
32'hBC199679,
32'hBE7CE5C1,
32'h3EA316B1,
32'h3D74D5FD,
32'hBED6B702,
32'hBD0DB376,
32'h3C990B1B,
32'h3F4F9161,
32'hBEFECDD8,
32'hBDD57F5E,
32'hBF4873AC,
32'hBD4CC625,
32'hBDA259F0,
32'hBE567C55,
32'hBD44EAA2,
32'hBD8C2710,
32'h3E7A27AB,
32'hBCD2F216,
32'hBD8ED63D,
32'h3D9997D6,
32'hBD7F43F1,
32'h3CF9A9CF,
32'h3CA2938C,
32'h3F388605,
32'hBE3D889C,
32'hBE041E27,
32'hBEBD1250,
32'hBEE46EEB,
32'hBE3473B3,
32'hBD04F827,
32'hBD8E7562,
32'hBE91119F,
32'hBCB403AA,
32'h3D6868AC,
32'h3E9A4838,
32'hBD562071,
32'h3D745214,
32'hBE23B0F3,
32'hBD9AF209,
32'hBD0C7E63,
32'hBDD7D4AF,
32'h3DC84924,
32'hBDA7AF1A,
32'hBD8F6A18,
32'h3CDC9AE0,
32'hBD506140,
32'hBD861A90,
32'h3C9CE572,
32'h3D9D9CD5,
32'hBD85BFC3,
32'h3D24C128,
32'h3C0CA7FF,
32'h3D2C5C2A,
32'hBD471EE2,
32'hBDAA5C82,
32'h3D84C1D3,
32'h1DDFB639,
32'hBC9A2E62,
32'h3D52B0BC,
32'h5DDD2957,
32'h1DC13A72,
32'h3D9084B5,
32'hBD461EEA,
32'h0EC1571A,
32'hBD5C0583,
32'h3D8E4C6E,
32'hBD87577F,
32'hBD292AAA,
32'hBDA73A60,
32'h3D29E4CB,
32'hBCD61907,
32'h1753070D,
32'h5DCC717D,
32'h3D237DAE,
32'h3DA45937,
32'h3C4861E4,
32'h3DD0FCBC,
32'hBD754C95,
32'h3D602369,
32'hBDD30219,
32'hBD5B840B,
32'h3DE0798B,
32'h175AE00F,
32'hBC3928FF,
32'hBD74826C,
32'h3D0AAF43,
32'h3DBD1FC6,
32'h3DA26AB7,
32'hBC9C6F4A,
32'h3D617031,
32'hBDB5CE45,
32'h3C9CF35C,
32'hBD9B2211,
32'h3DB37E02,
32'hBDDE84B5,
32'hBD1980D7,
32'h3D9C6656,
32'hBCC00FF5,
32'h3CD12919,
32'hBD301846,
32'hBD0827EE,
32'h3EE2953D,
32'hBDE1421F,
32'h3EF51271,
32'hBE29C144,
32'h3C902C2E,
32'h3CCA9E38,
32'h3E90CD26,
32'h3E83864C,
32'hBDC08B85,
32'h3F4FF8E5,
32'h3CE9C427,
32'hBD178243,
32'hBE939738,
32'h3F468C8F,
32'h3ED73665,
32'h3F696519,
32'h3E39776F,
32'hBDBE05C0,
32'h3C8172C3,
32'h3CB8835D,
32'hBE8AF1B7,
32'hBE0455E3,
32'hBF38D9B1,
32'hBF7B8F91,
32'h3EDDD945,
32'hBD50399A,
32'h3E5E49BC,
32'hBD7B50C6,
32'hBC18595E,
32'hBED96433,
32'h3F4A96B3,
32'hBE58102A,
32'hBE9E2A20,
32'h3E5BF665,
32'h3E629DD5,
32'h3CC4035D,
32'h3F16309F,
32'h3E751035,
32'hBE791DD9,
32'h3F1AAE79,
32'h3CA12024,
32'h3D9E422D,
32'h3E2CEEC0,
32'h3E10D84C,
32'h3D9B0C93,
32'hBD8E6FEE,
32'h3E99B559,
32'h3CEE8D41,
32'h3E6D7598,
32'h1DFAB29C,
32'hBE55C054,
32'h3C62527B,
32'hBF1DB886,
32'hBE6F7319,
32'h3F6C4551,
32'h3F17397D,
32'h3F7467D0,
32'h3E02F0D7,
32'hBE7D474D,
32'hBF5F07BA,
32'hBD8FE5BC,
32'hBECCA205,
32'h3F22F188,
32'h3F4C3E6C,
32'h3ED4C942,
32'hBF04FDA1,
32'h3F842356,
32'h3EDCEE04,
32'h3D405751,
32'hBF5BF1D8,
32'hBDB9F79E,
32'h5DDEE9FB,
32'hBF62B3A4,
32'h3F0D6CF3,
32'h3EE7C058,
32'hBEF78D26,
32'h3EC32E76,
32'h3E062DA3,
32'hBFBA26C4,
32'h3E1F9248,
32'hBD2E72EB,
32'h3E6ED209,
32'hBDBFB5BD,
32'h3EF10CCD,
32'hBD10F13C,
32'hBEC6F796,
32'h3DEA57AB,
32'h3F2F53BE,
32'h1DDA07EC,
32'hBC67127D,
32'h3E911A75,
32'hBF141D46,
32'hBF8CB376,
32'hBF4564BA,
32'h3DADDD10,
32'hBFAB6E46,
32'h3F5A8BE8,
32'hBED2B23E,
32'hBE5F176F,
32'h3E7D09CD,
32'h3D700A72,
32'hBD587812,
32'hBF08DCBF,
32'hBF047F07,
32'h3E947455,
32'h3E5220C6,
32'hBED01E01,
32'h3E14C7CD,
32'hBF10AE68,
32'h3D96B508,
32'hBEA72DE1,
32'h3E802A5E,
32'hBF248FC8,
32'h3E58DE79,
32'hBEA25EF1,
32'h3D8300A8,
32'hBEA7CA98,
32'h3ECB6535,
32'hBE956391,
32'hBE6877A0,
32'hBE8BC00D,
32'hBFBE54C5,
32'hBF184BBE,
32'hBE33C962,
32'h3E8A84D9,
32'hBF8C2E2B,
32'h3F04F760,
32'h3D31966A,
32'h3EB766FA,
32'h3EA4CDEF,
32'h17526F1F,
32'hBD0A8D2F,
32'h3EB61946,
32'h3E98B252,
32'h3DB6201B,
32'hBDA33E0E,
32'hBE2BFA97,
32'h3DC41A2C,
32'hBF81C8C2,
32'h3E25C05E,
32'h3D7DECE7,
32'h3EDCAECE,
32'hBF8BFC15,
32'h3E2870A2,
32'hBEC98EB3,
32'hBF178B49,
32'hBF19D0CA,
32'h3E38A3A6,
32'h3D871E3C,
32'hBF587907,
32'hBE53E197,
32'hBFB9B4E6,
32'h3ED04515,
32'hBE6E1C4E,
32'h3F3D2F51,
32'hBE1C44C0,
32'h3E5DF565,
32'h3E1CCF01,
32'h3E891D76,
32'hBE145D45,
32'h3A2814E,
32'h3DAE6D7B,
32'h3CF1EA13,
32'h3E8B6FA3,
32'hBE978F23,
32'hBE92E884,
32'h3EC93E1C,
32'h3CC81C7E,
32'h3DC6AE7E,
32'hBCEA3516,
32'h3EF4AF77,
32'h3E6B8E85,
32'hBFBE393F,
32'h3F086F44,
32'hBD9E8462,
32'h3D5518B3,
32'hBF22EF9C,
32'hBDF88A74,
32'hBE38297C,
32'hBF3DD70C,
32'hBFC459DF,
32'hBDCD63BF,
32'h3E4CF8C8,
32'hBE4BCF60,
32'h3F868EB4,
32'hBC674040,
32'h3CB25E46,
32'h3DB94F11,
32'hBE035260,
32'hBF46EA09,
32'h3D716CBF,
32'hBD6C35EF,
32'hBD272F4E,
32'hBC5894BF,
32'hBEDA164B,
32'hBDFAD68C,
32'h3D9CBF95,
32'hBEF2C79E,
32'h3F0B45F1,
32'hBE7ABFAD,
32'h3E5FEB84,
32'h3EF4F995,
32'h3F34ED8E,
32'h3E34C783,
32'hBE3F071A,
32'h3F51F565,
32'hBE2A5F0F,
32'h3D0F32A0,
32'hBE857433,
32'hBF00A7FE,
32'h3DB5EBF5,
32'hBDAA13D8,
32'h3E8966B2,
32'hBE645B43,
32'h3F3A2C30,
32'hBE4C66D8,
32'hBDE269ED,
32'h3ECB7D98,
32'hBEAFA959,
32'hBF153495,
32'hBD56C0FC,
32'h3D952EC2,
32'h3DF1E14E,
32'h3E77D5E9,
32'hBF21C742,
32'hBDFD9FD1,
32'h3E13B151,
32'hBDD23C07,
32'hBEB3DD53,
32'h3DC3A14F,
32'hBE81FED1,
32'h3E817849,
32'h3E81DCEA,
32'h3E6860DE,
32'hBE900F12,
32'h3EF207A6,
32'h3CA4E41D,
32'hBEF33E74,
32'h3DB916D2,
32'hBEC01A91,
32'hBFD987AB,
32'hBFA1398D,
32'h3E35ED33,
32'hBE3C4C22,
32'h3EA3F24A,
32'h3EE7ECF1,
32'h3D1039AE,
32'h3E47476C,
32'hBE2E54E8,
32'hBEF4F2F8,
32'hBD903819,
32'hBD3E41A4,
32'h3EB9F0DE,
32'h3E63D5AD,
32'hBE912D78,
32'hBDA783E6,
32'hBEC3EBC3,
32'h3E5C224D,
32'hBE8CA656,
32'h3C94437C,
32'hBE25B539,
32'hBD5D71ED,
32'hBDF3096C,
32'hBE8B674E,
32'hBE91A3C8,
32'hBEB4B51D,
32'hBE64973C,
32'hBCAC4985,
32'h3E240004,
32'hBE3EA7DC,
32'hBFD899C1,
32'hBE6C19C6,
32'hBC83BE6F,
32'hBE46ED95,
32'hBE301679,
32'h3D8728B3,
32'h3DD2F21E,
32'h3D80B3FB,
32'h3E806C0C,
32'hBD8CF343,
32'hBCC1B339,
32'h3CFCD1AF,
32'hBE58D396,
32'h3E0CA113,
32'hBEA541ED,
32'h3DB65696,
32'h3DB76BC4,
32'hBC710E08,
32'hBD119C40,
32'hBDAD0B72,
32'hBD6B4E7F,
32'h3D9F7087,
32'hBE4C2FB7,
32'hBD99178F,
32'h3D8655F6,
32'hBE633148,
32'h3E3CF3CE,
32'hBDAABA1B,
32'h3E510EA1,
32'hBEBDFEE6,
32'hBF6D6871,
32'h3C347932,
32'h3E7B8C4A,
32'hBCD37DA1,
32'h3DFEC402,
32'hBD43E353,
32'h3DC538C8,
32'h3EE86241,
32'h3E5DB390,
32'hBDADF3EB,
32'h3C80E3DE,
32'hBD0F8DD1,
32'h3D993244,
32'h3E5BA4B3,
32'hBE7C5956,
32'hBDD3520D,
32'h3E8C3C8A,
32'hBC917B17,
32'h3E3F84CE,
32'hBE9E49D2,
32'h3D3DC34D,
32'hBCCB6A35,
32'hBDAFFF95,
32'h3DEF5926,
32'hBE534E99,
32'h3DF2B922,
32'hBDA548B2,
32'hBE217E3D,
32'h3D1A9303,
32'hBF450CBE,
32'hBF808CEA,
32'hBF10CD7B,
32'h3DF4074A,
32'hBD51512D,
32'hBDC109D4,
32'hBDABAE92,
32'h3E665EC2,
32'h3EA2DDD5,
32'h5DCE0949,
32'hBE6CDD72,
32'h3D77C834,
32'hBDB3F47B,
32'h3E6C7640,
32'h3EAEC458,
32'hBE171E6A,
32'hBDE2B44E,
32'h3E603180,
32'hBDECF52F,
32'hBEB3EB97,
32'hBEA34AEB,
32'h3E30E489,
32'hBE15BDC2,
32'hBE92DE2D,
32'h3E359BD7,
32'h3C3028E8,
32'hBEDC41F1,
32'hBE7D0166,
32'hBE08F099,
32'h3D4FF6B1,
32'hBEC78978,
32'hBED88D35,
32'hBE99924A,
32'hBE3B8128,
32'h3CCE901F,
32'hBD2348C2,
32'h1751B18E,
32'hBD87DD5A,
32'h3DC7918C,
32'hBEC9B186,
32'hBD8B07EE,
32'hBDCA8B7F,
32'h3C9815DE,
32'hBE2A2FF2,
32'h3E99C743,
32'hBEAAF182,
32'h3D5010DF,
32'hBDBC1455,
32'hBF90155C,
32'hBE813648,
32'h3DFF1EC8,
32'hBD24B4FE,
32'hBCD55CC7,
32'hBE781EF8,
32'h3DAA9FA7,
32'hBDA88A9F,
32'hBEE83E89,
32'hBCF1AFFC,
32'hBCED0132,
32'h3E9892BE,
32'h3E6E5426,
32'h3E8B3646,
32'hBF6E9B30,
32'hBD85694C,
32'h3D8893AE,
32'hBE402689,
32'hBD819004,
32'h3E35D237,
32'h3E8A4E41,
32'hBE9F3B56,
32'h3E7671B0,
32'hBE19966F,
32'h5DC26AAE,
32'hBF000E33,
32'h3E79954D,
32'hBEAC9EBF,
32'hBCF6B99A,
32'hBED5FE6B,
32'hBF5526E5,
32'hBD7247F7,
32'hBE724DE6,
32'hBEAA24D8,
32'hBD76106A,
32'hBE9FA8FD,
32'h3C3629F2,
32'hBD8E1446,
32'hBE8BF07E,
32'hBEB16445,
32'hBF04247C,
32'h3E099594,
32'h3E60EA51,
32'hBDFC5013,
32'hBF2E30F5,
32'h3E056708,
32'h3E2EEA98,
32'hBF079BE1,
32'h5DCF499F,
32'hBD535270,
32'h3E8269F7,
32'hBCFA491E,
32'h3E6C4C64,
32'h3D3D71E0,
32'h2EC1B530,
32'hBF004B1D,
32'h3E9B318F,
32'h3E36DB32,
32'hBDBC3112,
32'hBE7B4AB5,
32'h3E88CD91,
32'hBE34EB46,
32'hBDAAA994,
32'h3EC87AA4,
32'h3E312451,
32'hBF0E4B52,
32'h3D5FCD65,
32'hBE2B470A,
32'hBF28C0F5,
32'h3E0B7494,
32'hBE370247,
32'h3E2D7F68,
32'hBEAD3F16,
32'hBDFC206B,
32'hBF8C23F0,
32'hBE2DD185,
32'h3D176952,
32'hBF26D526,
32'h3E26A623,
32'hBE06B52C,
32'hBE491E7A,
32'hBE2928A2,
32'hBDA2AB90,
32'h1DD03210,
32'h0ED85797,
32'h3D8C5C42,
32'h3D528F0F,
32'h3E0C1F3A,
32'hBE287C91,
32'hBE836FFA,
32'h3EC97595,
32'hBF23FE88,
32'h3E7CB7A5,
32'h3EADC390,
32'h3E7C844B,
32'hBD78B59B,
32'hBC847689,
32'hBD9DFCCE,
32'hBF145CEC,
32'h3E7B748A,
32'hBE62E77A,
32'hBDC2B9EB,
32'hBD877AD6,
32'h3C775803,
32'hBFC7123B,
32'hBE46023B,
32'h3C232C43,
32'hBEBB2C3A,
32'h3D987EF4,
32'hBC6BC8E4,
32'h3E17F0CB,
32'h3E13886C,
32'hBED703F3,
32'hBD3DF73B,
32'hBCE18BFB,
32'hBDC1052F,
32'h3D08A4F3,
32'h3E397344,
32'hBD526588,
32'h3E82DBBC,
32'h3E08896F,
32'hBE8ED740,
32'h3E9F863D,
32'hBF06044A,
32'hBE6FC71A,
32'h5DE4FAEF,
32'hBDF06A6D,
32'hBDF122CE,
32'hBF4C9160,
32'h3E6AC0A9,
32'hBF014C4E,
32'h3D9C6110,
32'h3E2A896E,
32'h3E248DE9,
32'hBF904243,
32'hBE3C48E0,
32'h3E9AB2B4,
32'hBDBFF239,
32'h3E38DF0C,
32'hBCB60D6F,
32'h3E3B68AE,
32'h3EDF7286,
32'hBEC4B0DD,
32'hBD6CDEF3,
32'h3D8514E3,
32'h1DCE043B,
32'h3EA0E282,
32'h3E8972EB,
32'hBE3D5B20,
32'h3D1F3FBD,
32'h3E33655B,
32'hBD60D031,
32'h3ED37AC2,
32'hBEA1CC51,
32'hBEA977E3,
32'h3C3F735D,
32'hBD04B5AC,
32'hBEB1036A,
32'hBFEDE605,
32'h3E4A8F46,
32'hBF2ECCE5,
32'h3EDB9E38,
32'h3E76C90C,
32'hBCAB931E,
32'hBF7B4681,
32'hBE6C744A,
32'h1DDFF9B8,
32'hBDA88FEE,
32'h3E11D173,
32'h3CEE8FD9,
32'hBDD8FE8A,
32'h3EAC8E38,
32'hBFD9C407,
32'hBD4F5CAE,
32'hBDD7A028,
32'hBDAED6B9,
32'h3E3E9B59,
32'h3E9EC0C4,
32'hBE4A2192,
32'h3EC2C787,
32'h3E7300F9,
32'hBEF57EB8,
32'h5DCD2EA5,
32'hBE455C37,
32'hBD3B1214,
32'h3F1260A8,
32'hBDBA92C1,
32'h3CC01AE1,
32'hBF63EF9A,
32'h3ECFBDB5,
32'hBEE12DF2,
32'hBE353247,
32'hBE951A25,
32'h3E22BF5F,
32'hBE8A8516,
32'hBE88B2A7,
32'hBC5E0074,
32'h2EC10C69,
32'h3E2627F5,
32'hBEA4060E,
32'hBD924E82,
32'hBEFC12B2,
32'hBFB61146,
32'h3D1F6E48,
32'hBDCCE050,
32'hBE8BC6EF,
32'h3EB64C59,
32'hBD5F3D33,
32'hBD59F4A5,
32'h3E65649E,
32'h3EA291B4,
32'hBED4C54F,
32'h3E42FE7A,
32'h3E228BF7,
32'hBCAECAAE,
32'h3D8D4310,
32'hBDD6C4CC,
32'hBF138E4F,
32'hBF7D59E3,
32'h3EF9AE7F,
32'hBE90A469,
32'h3E82A2E0,
32'hBD008709,
32'h3F413BF6,
32'hBF3C52ED,
32'h3D5A240B,
32'h3E1896A4,
32'hBCE3CA56,
32'h3EC0546B,
32'hBF1D604F,
32'h5DF2613C,
32'hBF67A6F7,
32'hBE826A29,
32'h3DAD29A5,
32'h3CFB6E33,
32'hBEC2FFF9,
32'h3E9B9C42,
32'h3EE1BBA3,
32'hBDB23BA5,
32'h3C4EB73D,
32'hBC62E441,
32'hBF567B2F,
32'h3ED3760D,
32'h3D96EAC5,
32'hBDBDBC2E,
32'hBE562EF4,
32'hBDF02D9E,
32'hBE985C2C,
32'h3E33FEE2,
32'h3F08F5DF,
32'hBC763BD3,
32'h3E1CC3BA,
32'h3C085BF2,
32'h3E801D73,
32'hBDB1B6A5,
32'h3F12F431,
32'h3DA33894,
32'hBE59731D,
32'h3F20E664,
32'hBF251BDE,
32'hBE7CBC0B,
32'hBFC16896,
32'hBEC60BC8,
32'h3D80363E,
32'h3D87F828,
32'hBEDF3A9E,
32'h3D121820,
32'h3E2A47EC,
32'hBE65C7CA,
32'hBD7FD136,
32'hBE034E96,
32'hBE65B655,
32'h3F332826,
32'h3EC82BD3,
32'hBE9D1265,
32'hBE9192B5,
32'hBEAB9D1C,
32'hBE628E37,
32'hBEDA13ED,
32'h3EB302D2,
32'h3DE7BEB8,
32'hBF23A57A,
32'h3EF33787,
32'h3E0296F9,
32'h3E70F9C8,
32'hBED14D7E,
32'hBEB43CFB,
32'h3E1E9E3F,
32'h3EE82F68,
32'hBF253D77,
32'hBF044EF4,
32'hBF24D631,
32'h3E0C5192,
32'hBD8049BF,
32'h2ED23C07,
32'h0ED9C554,
32'hBF75D9D7,
32'hBED19678,
32'hBE80261B,
32'h3D535FC8,
32'hBE82B06E,
32'hBE075673,
32'h3E11B66A,
32'h3EA14E9E,
32'hBE6896AD,
32'hBEBB262C,
32'hBE782A41,
32'hBF96AF8E,
32'hBE456AE6,
32'h3D0F170D,
32'hBDBC9990,
32'hBF3B6B4C,
32'h3ED5C792,
32'hBEE5B615,
32'h3F5121C2,
32'hBDE10AA4,
32'hBFCC604B,
32'hBE448C35,
32'h3DA676EE,
32'h3E236E9E,
32'hBEE6090C,
32'h3F1F86DE,
32'hBD777C76,
32'hBD8E41C5,
32'h3D52F8AB,
32'hBF35C17D,
32'h3F65747C,
32'hBF015D03,
32'hBD2DB877,
32'hBEC1283F,
32'hBDD0BDC2,
32'h3EB65829,
32'h3F7F29D3,
32'h3E71A560,
32'hBE1867EE,
32'hBF432014,
32'hBEF626F1,
32'hBF72E970,
32'hBEA59D01,
32'hBE462E85,
32'h3F2515D0,
32'h3EDCF703,
32'hBF0C03DA,
32'hBE47088B,
32'h3F16CA83,
32'hBF0679A3,
32'hBFBBA139,
32'h3E90CDDD,
32'h3F207F61,
32'h3D59E1BC,
32'h3F1A90A6,
32'hBD43E4FC,
32'hBD2DBF8D,
32'hBC1ED824,
32'hBD676DE9,
32'h3E95944A,
32'hBDE16601,
32'hBDA9193E,
32'hBF58BB0F,
32'hBF1D1796,
32'hBED7249B,
32'h3F11D054,
32'h3EB7D102,
32'hBFBFA446,
32'h3EE69796,
32'hBF203F06,
32'h3C520060,
32'hBD924613,
32'hBE5B4E30,
32'h3F3A05BA,
32'h3F5EB186,
32'hBD9B5486,
32'hBF2BDC0F,
32'hBDC8FFBE,
32'h3EA5391F,
32'hBE54EECE,
32'hBF41EBD7,
32'h2EC279A0,
32'h3E2EE5EA,
32'h3DE0914B,
32'h3E8863C2,
32'h3C15F021,
32'h3CF21276,
32'hBCA23AED,
32'h3C7D70B0,
32'h3F45B752,
32'hBE49166B,
32'hBDA05156,
32'hBF2AF90C,
32'hBF0633E0,
32'hBC18F6BF,
32'hBE50A167,
32'h3CAD14B8,
32'h3E3A0976,
32'h3DB3E35D,
32'h3E0EE508,
32'h3F30B609,
32'hBE364F78,
32'hBCD7794D,
32'hBECBFF8F,
32'h3EACF810,
32'h3D5FE8AB,
32'h3EBD660D,
32'hBCBCCCAC,
32'hBDC72182,
32'hBD65CD0A,
32'hBDBD9C65,
32'h3D23D6C7,
32'h3C8458B2,
32'hBD92F500,
32'hBD962E09,
32'h3DC02FE6,
32'hBC947D24,
32'h3D862AA0,
32'hBCDA2C6C,
32'hBC5D3243,
32'h2ED1D579,
32'h3DD7A1D1,
32'h2EC8D47E,
32'h2ED85A27,
32'hBC844CE2,
32'h3C884B72,
32'hBD9350DD,
32'h3D30798B,
32'h5DCE0C16,
32'hBD1E79DB,
32'h3D12F812,
32'h3CBF7642,
32'h3DA6C3DD,
32'hBD5F1A4C,
32'hBD4FD362,
32'h3C36554A,
32'h2EDB7542,
32'h3C813748,
32'h3C0CF323,
32'h3D28EB7E,
32'h3DE04434,
32'hBC94B116,
32'h175CA69A,
32'h3D92B9F2,
32'h3DD1A988,
32'h3D06DE23,
32'h3D31D1C9,
32'h3D264C0B,
32'hBDC5D2EB,
32'h3D6C44C7,
32'h3C248C29,
32'h5DE0494E,
32'h3CA977AB,
32'h3C79D844,
32'h3D9C6BDE,
32'h3CF89EFF,
32'h1DFC2EDF,
32'hBE348CA1,
32'h3E297CB2,
32'h0ED25039,
32'hBF200111,
32'h3F15EF39,
32'hBD0251B0,
32'h3EF01834,
32'h3D0E84EE,
32'h3D47A0A5,
32'hBC8E5A72,
32'hBDBC53F6,
32'h3D9C5AA5,
32'h1DEEC467,
32'hBEF87E8F,
32'h3DCF08D1,
32'h3F104EB8,
32'h3F9B2AE9,
32'h3E7EE29A,
32'h3C0382FE,
32'h3EC04BDB,
32'h3D1F31D9,
32'h3C88BB30,
32'hBF0C4F5E,
32'h3E5653D9,
32'h3F092EFF,
32'hBEBE9C7E,
32'h3E43CA5A,
32'hBE1D3834,
32'h3EB6803D,
32'h3ECE8877,
32'h1DEDDDB1,
32'hBDA1E4FB,
32'hBDA07163,
32'hBED42445,
32'h3F269678,
32'h3EB82CF3,
32'h3E092112,
32'h3E98AB5C,
32'h3EFC1B31,
32'hBDD0BF10,
32'h3F0802E7,
32'h3F20B9F8,
32'hBF577D5D,
32'hBF7310A3,
32'h3ED46DF6,
32'h3E6DA7CC,
32'h3F1DAEEC,
32'h3EE051E4,
32'hBEB2AF63,
32'hBE47FCA7,
32'h3DBA67A9,
32'h3D55BC4A,
32'hBE5520A3,
32'hBF1669EE,
32'hBF404F10,
32'h3E0872B2,
32'h3EAF027C,
32'h3E55F182,
32'h3FAD3C8E,
32'h3F175D91,
32'hBE6F297E,
32'h3ED778B6,
32'hBE1C0A84,
32'hBDB168CC,
32'h3DDC3985,
32'h3FAD5576,
32'h3EA37FDE,
32'h3EEB0150,
32'h3EC439D0,
32'hBEAB9B73,
32'h3F0B45CC,
32'h3F192F89,
32'h3D1C6C09,
32'h3EBD4847,
32'h3EBCFA23,
32'hBED48BB4,
32'h3ECBB968,
32'h3F656F7A,
32'h3EE3FAD1,
32'hBD37A0E5,
32'h3CB17EAF,
32'h3CB82F85,
32'hBF3831E0,
32'h3F0239E3,
32'hBE62418A,
32'hBF56F44F,
32'h3F29F7D5,
32'hBEFCE43B,
32'hBEFA7BCE,
32'h3E2E0E01,
32'h3E1B27AF,
32'h3E96514B,
32'hBE1AAB32,
32'h3D7B140E,
32'hBE8307DB,
32'h3F21526A,
32'h3E3D6C21,
32'h3DB6F4AF,
32'h3DF5345E,
32'h3D52543D,
32'h1DCB1584,
32'h3F14AA1A,
32'hBE656701,
32'h3E11CA6B,
32'hBD777092,
32'hBF96E937,
32'h3F0DD698,
32'hBE178E71,
32'hBDE78F3C,
32'hBF2C7C6F,
32'h3DB4B79B,
32'h5DEBDFB2,
32'hBEB8C36A,
32'h3E106624,
32'hBE546CB5,
32'hBE8E0738,
32'hBEC38481,
32'h3E94FD5E,
32'hBE44D601,
32'h3EC9AF3C,
32'h3F459F46,
32'h3E69870A,
32'hBF808D09,
32'hBD44075A,
32'hBE84A015,
32'h3F78B563,
32'hBED423C6,
32'hBCC81A94,
32'hBDBE08B5,
32'h3EE084B7,
32'hBF15F621,
32'hBE11EF0E,
32'h3D82F59B,
32'hBDABF4D7,
32'h3E28D75F,
32'hBE422B80,
32'h3EAD939B,
32'hBEC24CFE,
32'h3E33FAAF,
32'hBEBBBC0D,
32'h2ECC2A8A,
32'h3C98D183,
32'h3CBF5332,
32'h3DF59A9A,
32'hBEB9EF3B,
32'hBD82ADFD,
32'hBCF20B3B,
32'h3E0F6173,
32'h3E6EC1B9,
32'h3C5AAF09,
32'hBD5FB5AC,
32'h3E6FA466,
32'hBF931AAB,
32'hBE8E1926,
32'hBDF385B7,
32'h3EABEBC8,
32'hBEF4AAF5,
32'hBECCEFBE,
32'h3EDF9F9A,
32'h3D3704F4,
32'h3D68B505,
32'h3C25C30F,
32'h3D063D6A,
32'h3DB80DD1,
32'h3EE61BBD,
32'hBF3703E3,
32'h3EAD03D7,
32'hBCDD7DAE,
32'h3E8418B1,
32'hBF58404C,
32'hBC84D43C,
32'h3C4DFA7F,
32'h3D0A2609,
32'hBE0DCD8F,
32'hBF0400F1,
32'hBE3263AF,
32'h3CEEFD29,
32'h3C789722,
32'h3EBCF715,
32'hBD9BFACF,
32'h3C2FD47C,
32'hBD731542,
32'hBF00CD77,
32'h3E8B2748,
32'h3D0A776A,
32'h3E69897B,
32'hBD236769,
32'hBF1B0898,
32'h3E2DA8F4,
32'h3D162E04,
32'hBEC2BF89,
32'h3A0FF81,
32'h3E334B57,
32'hBE33D3AA,
32'h3ED34710,
32'hBEB911D1,
32'h3E508816,
32'h3E357600,
32'hBD5A53E5,
32'hBEBC4C25,
32'h3DB64267,
32'hBCFCF006,
32'h3DE21ECF,
32'h3D28B6DA,
32'hBDCDA700,
32'hBD535276,
32'h3E8902DC,
32'h3D93D1DD,
32'hBCD1D18F,
32'h3E69CC01,
32'hBE942F6A,
32'h3E850CF3,
32'h3DA39FE5,
32'hBD7E8F09,
32'hBE2ED8EF,
32'h3E8029E7,
32'h3EAB801E,
32'hBF3EC9F4,
32'hBEA2992D,
32'hBEB56C97,
32'h3ED77139,
32'hBF502DF1,
32'h3EAE6E57,
32'hBF062ED2,
32'h3DB307B9,
32'hBEDBE523,
32'h3E86C260,
32'hBDA5D27A,
32'h3D2AED05,
32'hBEED5B97,
32'hBDCAFDCE,
32'hBCA304EA,
32'hBE5BBCEC,
32'h3D43B92F,
32'hBD2B0915,
32'hBDBE3463,
32'h3DFDC87A,
32'h3EBFEC46,
32'h3DDA310B,
32'h3E41429A,
32'h3E665833,
32'hBD412C9D,
32'h3EA27851,
32'hBE676811,
32'h3E846BBC,
32'h3EDD5FEA,
32'hBD79EDBF,
32'hBEC38827,
32'hBDDADFD5,
32'hBE674A0B,
32'h3E8A9CE9,
32'hBF1D3916,
32'h3D794F01,
32'hBDAB92CA,
32'h3DAC14E1,
32'h3D251D87,
32'h3D174FC4,
32'h3EA15F50,
32'h3E003621,
32'hBF69745F,
32'hBC9A6C60,
32'h3D4AC16F,
32'hBDEAC50F,
32'hBE0528FA,
32'hBE2D8055,
32'h3E53612E,
32'hBDFFCD60,
32'hBE956F20,
32'hBE44B2B6,
32'hBD61282A,
32'hBEDB4338,
32'h3EAE44AC,
32'h3E14BBF7,
32'h3D310DFF,
32'h3E0D450A,
32'hBDCF262F,
32'h3E66ABA5,
32'hBE082C67,
32'hBE216448,
32'hBF2C6626,
32'h3E6F1797,
32'h3D0DC135,
32'h3D70BC7B,
32'h3C9C0AE5,
32'h3ECD55C6,
32'h3E851AC4,
32'h3E1574D0,
32'h3DA2E969,
32'h3EF4D105,
32'hBE5669A5,
32'hBD2210EA,
32'hBD2D76BB,
32'h3CA2C501,
32'h3E34640E,
32'h5DED8DBD,
32'h3E6843E1,
32'hBEA6425B,
32'hBE433DC1,
32'h3DA30CDF,
32'hBDD41724,
32'hBF2CC7F3,
32'h3CB0B7BF,
32'hBE36BDE4,
32'hBDEEE0E9,
32'h3CD7FC41,
32'h3E37F267,
32'hBC32674B,
32'hBE23ECF4,
32'hBE2F7023,
32'hBF24FEC6,
32'hBF6DC8A2,
32'h3DB79226,
32'h3DF2FFD3,
32'h3C7D24FF,
32'h3EB04065,
32'hBDD60695,
32'h3DDC25ED,
32'h3E85BAD4,
32'h3E6DCF50,
32'hBC96554A,
32'hBCA4C1C9,
32'hBD48E8F7,
32'hBCBB3105,
32'h0EC13448,
32'hBD96529C,
32'hBE0C969E,
32'hBD6A7D5A,
32'hBEB6A5EF,
32'h5DCB696E,
32'hBEB3DFB6,
32'hBE65FD5B,
32'h3D04597F,
32'hBCA78E83,
32'hBE310C5F,
32'hBE441D76,
32'h3ECDD18B,
32'h3CFE611B,
32'h3E36E66B,
32'h3E0FF011,
32'hBEC5E26D,
32'hBF95E1A1,
32'hBE098234,
32'h3D1558D2,
32'h3DB7316C,
32'h3D01F983,
32'hBE3D0058,
32'h3E71C147,
32'h3E4E9591,
32'h3E18050D,
32'hBE253B2E,
32'h17557A31,
32'hBD237F24,
32'h3D83800E,
32'h3E2923A9,
32'hBDD1210D,
32'hBE023698,
32'hBDA6CB61,
32'hBED2A29C,
32'hBD04EC48,
32'hBE2FDFCE,
32'hBE63E49F,
32'hBCA1EADB,
32'hBF13D8E9,
32'h3C4924EB,
32'hBD8E283E,
32'hBE826EEC,
32'h5DDC3E7F,
32'h3E624421,
32'h3D00B3C4,
32'hBEA4A2E2,
32'hBEA2DD66,
32'hBE2331EB,
32'h3D292673,
32'h3E8622BC,
32'h3CF66AB6,
32'hBD9F58FB,
32'h3E4E5C8D,
32'h3C4C8945,
32'h3D08A5E4,
32'hBDD4A5F0,
32'hBD965B18,
32'hBD5F0F42,
32'hBE86B23D,
32'h3E0D00F0,
32'hBE379410,
32'hBDEA4905,
32'hBE14D245,
32'hBF2E6C07,
32'h3DC87E4E,
32'h3E3535A4,
32'hBE09C640,
32'h3C854952,
32'hBD5A3019,
32'hBE81ABD5,
32'hBD9784AF,
32'hBF0E1CB3,
32'h3D6E3848,
32'h3DA08876,
32'hBDFB8D38,
32'hBF12BB29,
32'hBED2DE67,
32'hBE4B7DC3,
32'h3CB33246,
32'hBC419900,
32'hBE454605,
32'hBE95A335,
32'hBCF5F2CD,
32'h3C95F351,
32'hBE7C07A5,
32'h3D55F715,
32'hBC96CF7F,
32'h1DD5A707,
32'hBE994189,
32'h3E424B76,
32'hBDA78131,
32'hBD9BB15A,
32'hBE8A21AF,
32'hBFDE4DED,
32'hBD0D8BD7,
32'hBEE8CA7D,
32'hBE596471,
32'hBDD0F812,
32'hBE5EEEEB,
32'hBD9B008C,
32'h3D455392,
32'hBE23209F,
32'h3E5E58DE,
32'hBE929F7F,
32'h3E116B11,
32'hBEF822AB,
32'hBE28B3F6,
32'hBEB4A0DA,
32'h3E3DA5DA,
32'hBE367DB3,
32'hBE488681,
32'hBE060CF8,
32'hBE934224,
32'h3E9B129C,
32'hBDBEE854,
32'hBE866932,
32'hBD5D1E7E,
32'hBD9B5646,
32'hBEAE5772,
32'h3E0C3568,
32'h3CAE834B,
32'hBD9A9B11,
32'hBD8703A7,
32'hBE6F7184,
32'hBD76F92E,
32'hBEC33293,
32'h3D21D7A0,
32'h3E11CAB7,
32'hBF1DB6C2,
32'h3D17E9E1,
32'h3E1092E9,
32'hBD014ABD,
32'h3E5C3EE4,
32'hBEA905ED,
32'h3E546001,
32'hBEE9411A,
32'hBE1BD26E,
32'h3E7C30F5,
32'h3D6C4EB5,
32'hBD47E0DE,
32'hBA54A31,
32'h3E4C17FB,
32'hBD98BD42,
32'h3C9BBA59,
32'h3EBD5903,
32'hBED683E4,
32'h1DDCBF84,
32'hBDA250E6,
32'hBF0E7DD1,
32'h3D3EAA83,
32'h3DB424A2,
32'hBCB87A89,
32'h3DF2483A,
32'h3D86C598,
32'h3F0F10FF,
32'hBEB0BD18,
32'hBE1922EA,
32'h3E402DF4,
32'hBE286E03,
32'hBEA9E616,
32'hBDC1A7ED,
32'hBD456CAB,
32'h3E05B1F0,
32'hBDC698CF,
32'h3DA82763,
32'hBEE9D9E9,
32'hBE0329FC,
32'h3ECC28CC,
32'hBE084E16,
32'h3E08FBC8,
32'h3CFDBEEC,
32'h3E7256D2,
32'h3D05F36E,
32'h3CADFE71,
32'h3E1670B3,
32'hBDD8301F,
32'hBDB02838,
32'hBD0DFBE2,
32'hBE9994FC,
32'h3E6A70A7,
32'h3DB6AD18,
32'hBD220065,
32'h3EDEFC04,
32'h3DBCB526,
32'h3EACFA87,
32'hBEF833F7,
32'hBEFF9E72,
32'h3C1335C1,
32'h3DE07422,
32'hBEBD1630,
32'h3E5B8881,
32'hBE68ECF1,
32'h3E7DE9B2,
32'hBD8CF76B,
32'h3DDD8FD4,
32'hBEFBA76C,
32'hBC6E601C,
32'h3D1E69E1,
32'hBE124B39,
32'hBE9F13FD,
32'h3E6D4BE3,
32'h3E3E248B,
32'hBE12D9D0,
32'h3E325820,
32'h3EF259E1,
32'hBEF14AA3,
32'h1DC1E6BB,
32'hBDF71F92,
32'hBE232C8E,
32'hBDDC361F,
32'h3E62D3D5,
32'hBE96C6F3,
32'h3D91F129,
32'h3E3470A8,
32'hBE0FA264,
32'hBEDB99D5,
32'hBF1E1D30,
32'h5DEBE80C,
32'h3E6D81E3,
32'hBD8227BE,
32'hBCDA57D6,
32'hBD9C7C0C,
32'h3E560CDA,
32'h3D0FB638,
32'h3CFF2C48,
32'hBD828AA2,
32'hBE3A24EE,
32'hBE1CAD30,
32'hBF059C43,
32'hBEB73B53,
32'h3E3635E7,
32'h3D93030D,
32'hBD9D9052,
32'h3E3A6E96,
32'h3DC29B73,
32'hBFC6C356,
32'hBCFECCC5,
32'hBC80A160,
32'hBDE3E0CE,
32'hBE99CAE8,
32'h3E240AB8,
32'hBD95E81D,
32'h3DB12645,
32'h3DE7A56B,
32'hBE9BF17B,
32'h3C1C46BA,
32'h3DC8E0E8,
32'h3E3773FB,
32'h3EBCD839,
32'hBE33D1B2,
32'hBE147463,
32'hBE53EBFE,
32'h3E870B1A,
32'h3D897317,
32'hBE5AECF3,
32'hBE988838,
32'hBE415987,
32'h3E15E90C,
32'h3D57F61F,
32'hBC28B131,
32'hBDA65A9A,
32'h3E4A654B,
32'h3E649C8C,
32'hBCE2B2AE,
32'hBEB3B48A,
32'h3DAB6E1E,
32'hBDDC1FDD,
32'hBC6E585C,
32'h3C1F3A1C,
32'hBE93F0A4,
32'h3E26ED1A,
32'hBC82F7D0,
32'hBD188295,
32'hBD51C45E,
32'h3E150917,
32'h3CF63D01,
32'hBE0123F0,
32'h3CDA09C1,
32'hBF34D3BB,
32'hBE51CF36,
32'hBEC1ABFD,
32'h3DAFA558,
32'h3E759E6F,
32'h3EA4C43D,
32'h3EB46402,
32'h3E0DF1F3,
32'h3D5F1FC4,
32'h3EAA5E25,
32'h3EC04218,
32'h3EC47813,
32'hBE334784,
32'h3DC66567,
32'hBE9B280D,
32'hBD2DD5DC,
32'hBF80E90F,
32'hBF325E38,
32'h3D614B02,
32'hBD08BAEB,
32'hBE8F6958,
32'h3E7E701E,
32'hBDF282BA,
32'hBE5102C8,
32'hBE893335,
32'h3E816704,
32'hBEC55B74,
32'h3CFA1869,
32'h3DC0888B,
32'hBD1CDEBA,
32'h3E3FBA9C,
32'hBE38C490,
32'hBE01D636,
32'hBF4D3251,
32'h3D6371EE,
32'h3EA0D489,
32'h3EBB25B2,
32'h3E87D9AC,
32'hBE83F7ED,
32'hBE430C39,
32'h3C288248,
32'h3E44A9AC,
32'h3DA08517,
32'h3EFB2A5D,
32'hBFC781AA,
32'hBE14DEE1,
32'hBFFA142C,
32'hBEF26E5E,
32'hBD982EB9,
32'h3DAFE2BD,
32'hBF719159,
32'hBF07BF28,
32'hBEE8D304,
32'hBDFDFDE9,
32'hBE19F039,
32'h3E8B43B8,
32'hBF71F741,
32'h3EBB8E17,
32'h3EF4A2B4,
32'h3CA48CFE,
32'hBD0295D1,
32'hBE0EC415,
32'hBEA92A68,
32'hBF090326,
32'h3E248329,
32'h3DA037EE,
32'hBF5B8969,
32'h3D7D12DA,
32'hBEFDAF76,
32'h3DCA92AC,
32'hBE5DA37D,
32'hBF0464A1,
32'h3D2AF1BB,
32'h3EB1D6C1,
32'hC0287CD8,
32'h3EC760EB,
32'hBFCD3541,
32'hBEBBFFBA,
32'hBDBBFCC1,
32'h3CAFD6AA,
32'hBFAC3AB5,
32'hC00DA289,
32'hBF78291C,
32'hBE4374B1,
32'h3E63AAB0,
32'hBF33CF41,
32'hBF04B867,
32'h3EAD1C6F,
32'h3EA0530F,
32'hBA28808,
32'hBD6E4188,
32'hBEA26D32,
32'hBF278E86,
32'hBCD24C15,
32'h3EBB3C1D,
32'h3E34EBE1,
32'hBF90D978,
32'hBF1B5922,
32'hBF14E102,
32'h3E911933,
32'hBFF26F7C,
32'hBFE5D6BC,
32'hBF9D1768,
32'h3F61B71F,
32'hBF8CC632,
32'hBD894F45,
32'hBECEAEBD,
32'h3EB69F16,
32'h3D3E2FDD,
32'h3D84580D,
32'hBF63683A,
32'hBE949C16,
32'hC0192FB8,
32'hBE3A493D,
32'hBF394F3D,
32'hBE846870,
32'hBD988D36,
32'h3E878BD6,
32'hBEDA9648,
32'h3E319FC1,
32'hBF4B9CF9,
32'h3E8E1FBD,
32'hBFA61925,
32'hBE9BF6D1,
32'h3F304973,
32'h3E00A785,
32'hBE984292,
32'hBF1A13A8,
32'hBF01091E,
32'hBF1D19FE,
32'hBDD480A8,
32'hBFC5FB61,
32'h3E53B4DF,
32'h3F776CF5,
32'hBE0FCA89,
32'h3E1731F4,
32'h3C2EB0CA,
32'h3E5CB3B3,
32'h1759224B,
32'h3D79075D,
32'h3F25D0C9,
32'h3E1B153D,
32'hBE870401,
32'h3E7D1FE8,
32'h2EC37333,
32'hBDCCEDB8,
32'hBEC448E0,
32'hBC662804,
32'h3FD1567F,
32'hBEB6F8E6,
32'hBF210FE9,
32'hBF5D012C,
32'hBEF2639E,
32'hBF0C575F,
32'h3EA1DA37,
32'h3EE61E9B,
32'hBD40D635,
32'hC0034476,
32'hBF0AC150,
32'hBED139A7,
32'h3E90B2E2,
32'hBF412502,
32'hBF6AF9B0,
32'h3DED9FEA,
32'h3D4BAE13,
32'hBEA5B5CC,
32'hBCA3FA88,
32'h3EC69EE5,
32'h3C863892,
32'h0ECFFEF0,
32'hBE44679C,
32'h3E3CFE75,
32'hBE36259E,
32'h3FA0B747,
32'h5DDB7293,
32'h3E895FA0,
32'hBF59CE83,
32'hBF967317,
32'h3F3E82AC,
32'h3FBA00D4,
32'hBE563197,
32'h3ED8DC7E,
32'hBEC0FDA5,
32'h3DAA817A,
32'h3E230C8E,
32'h3F73EBFA,
32'h3C352821,
32'hBF691703,
32'hBD8D9DA6,
32'hBC8B1AE6,
32'hBC82925C,
32'h3CEE90CC,
32'hBC07EE7E,
32'hBD0C700B,
32'hBD485F7D,
32'h3D9E6BF9,
32'h3DAE8F4F,
32'hBD09196E,
32'hBD1C62A3,
32'h5DCA1BAD,
32'h1DDE6A21,
32'h3D0EB773,
32'h3C1E015A,
32'h3C801AA1,
32'h0ED77545,
32'hBD4190E5,
32'h3D7AD106,
32'h3D1769AB,
32'hBDAC073D,
32'hBD9F85F6,
32'hBD22739D,
32'hBCBB0F37,
32'h3DB02441,
32'hBDC12CD9,
32'hBD0850FC,
32'hBCFEDCA5,
32'h3D039436,
32'h3D64D041,
32'hBCA9FA79,
32'h3EE64C19,
32'h3E7E5B01,
32'h3DB9EF0C,
32'h3EA6C185,
32'hBD8837BE,
32'h3FBF79EA,
32'h3FD7B4E7,
32'h3D50CC33,
32'hBD41DBFB,
32'h3CCA5029,
32'hBD6E4BC6,
32'hBF17D8D7,
32'h3DE4C4C0,
32'hBD4C6643,
32'hBFA65216,
32'hBD43F9DF,
32'hBDC3C777,
32'h3DD092E2,
32'h3E5CB8CF,
32'hBEEE0214,
32'h3E21E807,
32'hBD9FFB00,
32'hBFE85A3E,
32'h3FABDB79,
32'h3FD47F7F,
32'h3F0A77EE,
32'h3E84B274,
32'h3D126D00,
32'hBEF682A6,
32'h3D888332,
32'h3F1AC2EC,
32'hBDB03015,
32'hBF09F8DE,
32'h3EB4ADF1,
32'h3ED17CEB,
32'hBE675EBA,
32'h3E8715CC,
32'hBDD0E31D,
32'h3F2D031F,
32'h3C38DAC5,
32'h3DE6278B,
32'h3FBE14E8,
32'h40080846,
32'h3FBAB7B9,
32'hBF155307,
32'h3E0D6CFB,
32'hBE3A17FA,
32'h3ED45F68,
32'h3F3C723A,
32'h3DB1E974,
32'hBD9E0D43,
32'h3D5BE843,
32'hBF6B2D30,
32'hBE8E2977,
32'h3F628CF0,
32'hBE7092F6,
32'h3ED75C74,
32'h3F27F8F4,
32'hBED7528E,
32'h3F0D159E,
32'h3F736865,
32'h3F4ED0F9,
32'hBF17A91E,
32'h3F30393D,
32'h2EC424D1,
32'h3F370EC3,
32'h3F8613E7,
32'h3F22A44F,
32'h3EBF8985,
32'h3CCF80EC,
32'h1758CF04,
32'h3DA922AB,
32'hBF7ADC17,
32'hBEBCC80A,
32'hBE79DEAE,
32'hBF465626,
32'h3DC04F3C,
32'h3FA744C4,
32'h3CFA253F,
32'h3E054D3C,
32'h3E38B72C,
32'h5DC213F3,
32'hBF883D58,
32'hBF0ED944,
32'h400770FE,
32'h3EEBF8B1,
32'h3F198113,
32'h3EB76EC8,
32'hBE585E31,
32'h3F2472B5,
32'h3D8DE353,
32'h3DF79A74,
32'h3EECD957,
32'hBE8B17BB,
32'hBF67E915,
32'h3F0DB25D,
32'h3F0AD43D,
32'h3F09E122,
32'hBE17AC64,
32'h2ED00CFE,
32'h3D4F605D,
32'hBF8030F4,
32'h3ED041C5,
32'h3EC489CF,
32'h3E64086C,
32'hBEAB9E3B,
32'hBED15DCB,
32'hBEE35668,
32'hBD686842,
32'h3F0961A3,
32'h3E7A7A82,
32'hBE8E3516,
32'hBEC73B29,
32'hBF041ADF,
32'h3E3D3458,
32'h3F1EBE72,
32'h3D0EBBC7,
32'hBD36624C,
32'h3F4AEB84,
32'h3E096C6E,
32'hBE83C0A6,
32'hBA455F5,
32'h3EFCE525,
32'hBEEC1FBC,
32'hBF0A2644,
32'h3EB35438,
32'h3D92DC9F,
32'h3D8690BB,
32'hBF7DDB1C,
32'hBD904B28,
32'hBD727A58,
32'hBF1FA722,
32'hBE15BA53,
32'h3F15F89E,
32'hBE39C689,
32'hBEA92ECA,
32'h3E896DC4,
32'hBE2581DE,
32'h3E99D714,
32'h3ED63503,
32'h3EABD2CE,
32'hBF00CA3E,
32'hBD74BFF7,
32'hBE1DA1CF,
32'h3D30E05F,
32'hBE4BBB64,
32'hBF243FE3,
32'h3EB3F4C6,
32'h3E9582A2,
32'h3D3261C9,
32'h3E931C97,
32'h3DE81EA2,
32'h3E98A03D,
32'hBDB152CB,
32'hBC84EA5B,
32'hBD8DCD37,
32'hBECBD6A7,
32'h3E6475D8,
32'hBEC33C8F,
32'hBD315BA4,
32'hBC9283F5,
32'hBE36A3CD,
32'h3E94F335,
32'hBEBECCD9,
32'hBD5A4CFD,
32'hBE8CE05B,
32'h3EB10626,
32'h3F15DE38,
32'h3D8539CF,
32'hBE852E58,
32'h07590E76,
32'hBF8C9D13,
32'hBEAD0D1C,
32'h3D1DED17,
32'h3F0811D8,
32'hBE99948B,
32'hBE073352,
32'h3F456807,
32'hBD030DFD,
32'h3E12363B,
32'h3F68F5D8,
32'h3DB34B06,
32'h3E176A6B,
32'h3CCC41F4,
32'hBEFF49ED,
32'h3E151867,
32'hBEA973D8,
32'h3E650756,
32'h3E592255,
32'h3D895EBA,
32'h3D2CA199,
32'h2ED1BEFD,
32'h3E7D8CE4,
32'hBE60D8C1,
32'hBDC83CC0,
32'h3D1F44C4,
32'h3D375495,
32'h1DEFD754,
32'h3D5047CD,
32'hBF03DE0A,
32'hBC89BE63,
32'hBE55348C,
32'hBC8108D7,
32'hBD6FA6EA,
32'h3EC094F9,
32'hBE3CFB37,
32'h3F1C7618,
32'h3F0A768E,
32'hBD80D3EA,
32'h3DD67409,
32'h3E64A424,
32'hBE5F4346,
32'hBF02AA6B,
32'hBE902415,
32'hBEAA1FB4,
32'h3C81F635,
32'hBEDDB86F,
32'h3E04DDFB,
32'hBE1527C7,
32'hBD242CC8,
32'h3C416DAE,
32'hBE27EB5C,
32'h3E3D4C9F,
32'h3D09026A,
32'hBE0802D9,
32'h3E6D62A6,
32'h3DE713E9,
32'hBECCF09B,
32'h3E277698,
32'h3E3A5959,
32'h3D98A876,
32'hBEFF656F,
32'hBE25EB38,
32'h3DFD0D4E,
32'hBDBC7307,
32'h3EC9B88E,
32'h3D77892C,
32'h3EAA1D3A,
32'hBE91E1EC,
32'h3ECDC940,
32'hBD3732F6,
32'h3D8B1DFB,
32'hBE014224,
32'hBEA300EE,
32'h3DDBFE47,
32'h3D7BCCE5,
32'hBEB048C9,
32'hBC4A1F3F,
32'h3E4D3B64,
32'h2EC4CFCD,
32'hBD418591,
32'hBE881B5A,
32'h3E296F15,
32'h3E21D495,
32'hBE5F22B8,
32'hBD5AB74B,
32'hBE80D634,
32'hBDED90D4,
32'h3CC25904,
32'h3EBFB215,
32'hBE02FB9C,
32'hBD8F26F6,
32'hBE80A177,
32'h3EE86819,
32'h3F431852,
32'h3E08AD7C,
32'hBE595852,
32'h3E09EADE,
32'hBF5AD949,
32'hBE76BE98,
32'hBEAEA994,
32'h3D04CB6B,
32'h3EA24380,
32'h3D20D8BB,
32'h3EFEBEF5,
32'hBDDCC841,
32'hBD9F0A1C,
32'hBE915B82,
32'hBE364BF0,
32'hBD869A2C,
32'hBD8E2E41,
32'h3C18973C,
32'h3DDDF45B,
32'h3CC85890,
32'hBC124D26,
32'h0EC5A7B6,
32'h075B5F66,
32'h3DD9EF77,
32'hBE724E57,
32'hBE88118E,
32'hBDE073D4,
32'hBF423B89,
32'hBE22CB96,
32'hBD6E1EDF,
32'h3F06406A,
32'hBE65927D,
32'hBD972624,
32'h3CBEB9D7,
32'hBF34AD71,
32'hBE773FA9,
32'hBEC50AED,
32'hBDF6F9DF,
32'h3E8297D1,
32'h3EA97CEC,
32'h3E5CCCAD,
32'hBD9D3BF1,
32'hBF075A4A,
32'hBD4D8F8B,
32'h3C8452A3,
32'h5DD34DD6,
32'hBDADFD1A,
32'h3E624F19,
32'h3EC160F3,
32'h3DAB2735,
32'h3D775AE2,
32'h3C70E39A,
32'h3E147974,
32'h3D8A9583,
32'hBE2E38E3,
32'hBE9068F8,
32'hBDEB668B,
32'hBEECC097,
32'h3DF4A0FD,
32'h3EB25DC2,
32'h3E226D79,
32'hBE027EF6,
32'hBE3877D0,
32'h3D710F31,
32'hBF07C77A,
32'hBEAF2844,
32'hBF1187B9,
32'hBDED215D,
32'hBD92E6CF,
32'h3E3657CF,
32'h3DDBA4CD,
32'h3E15511D,
32'hBE5DFC06,
32'hBDA0B2AC,
32'h3EDA505D,
32'h3D94D3F0,
32'h175BF1E9,
32'hBE7735F7,
32'hBDAF4364,
32'h3D867D52,
32'h3DBB1292,
32'h3E37786D,
32'hBD7729C6,
32'h3E50C8A1,
32'hBECC7F9E,
32'hBF04C9C3,
32'h1DE8AFB2,
32'hBF1293D3,
32'hBDA49A16,
32'h3E15BF92,
32'hBE1E2C45,
32'h3D363F29,
32'h3E56B2B1,
32'hBE70F07C,
32'hBECE1CEE,
32'hBE8E0FF8,
32'hBEDCCB0E,
32'hBD5A224F,
32'h3C4BC56C,
32'h3E34279E,
32'hBE904047,
32'h3E8A43A3,
32'hBE37E44F,
32'h3E3AC4D9,
32'hBE72FA4D,
32'hBD9FF35F,
32'hBDA21708,
32'hBE26B068,
32'h3E91E337,
32'h3C39977F,
32'h2EC57CF6,
32'h3E107813,
32'hBD253D30,
32'h3E18FA63,
32'h3C982924,
32'h3C8E6BA6,
32'h3E589535,
32'hBEE59A58,
32'hBE05BD82,
32'h3E8ECA1C,
32'hBE765338,
32'hBD8A525A,
32'hBCAD193A,
32'hBE2DD66D,
32'h5DE81FE3,
32'h3C96B738,
32'hBE6E96CA,
32'h3D9E9071,
32'hBD8DF5B0,
32'hBE5362C1,
32'hBD6CEA5F,
32'h3E2F6008,
32'hBDA23CF1,
32'hBD3BE16B,
32'h3DC8B9E1,
32'h3CAA094C,
32'h3DA9AAAE,
32'hBE176CCF,
32'h3E2E96B1,
32'hBE579C44,
32'hBE9C8D3A,
32'hBD25C6D0,
32'hBF8E1A35,
32'h3E1E74CE,
32'hBE2AEADC,
32'hBE1DF718,
32'h3D6C51A6,
32'hBDDD30B4,
32'hBD19DFE8,
32'h3E713BAF,
32'hBEF55DA3,
32'h3C66981A,
32'hBEA13996,
32'hBD1AD535,
32'hBE9BCF13,
32'hBE8174BB,
32'hBE316B54,
32'h3D2C538B,
32'h3DC01C04,
32'hBE9D15FD,
32'hBEA02463,
32'hBEDCA664,
32'h3DED5A99,
32'hBE742ED1,
32'h3D2D9E42,
32'h3D3C01D3,
32'h5DDE0C4A,
32'hBE592A70,
32'h3E1122F0,
32'h3DB58859,
32'hBD0FFE51,
32'hBEE006C1,
32'hBF90F601,
32'h3C216F6F,
32'hBEB1C4D5,
32'hBC8BA0AC,
32'h3CA1D27F,
32'hBDF0A55F,
32'hBD1A0B19,
32'hBE011B60,
32'hBF0F1E88,
32'h3D6F08F8,
32'hBEFD2D9C,
32'h3D780029,
32'hBF07EEF5,
32'h3D909C00,
32'hBE33406E,
32'h3DDE7D79,
32'hBD02A61E,
32'hBE86516F,
32'h3D615C2B,
32'h3D87EF91,
32'h5DE0C6DC,
32'hBEE56232,
32'hBD33FC4A,
32'hBE09CAD8,
32'hBD8EDA3F,
32'hBF263D7D,
32'h3E2FBEEC,
32'hBE0CCDCC,
32'hBE1DFB9D,
32'hBDB8D340,
32'hBEEA5BCC,
32'h3E8F260D,
32'hBE9D6D69,
32'hBE095E8A,
32'hBDD95FD6,
32'hBF16E131,
32'hBE48E64B,
32'hBE00B273,
32'hBE838EF8,
32'hBD1E0429,
32'hBE436729,
32'h3E7AD366,
32'hBE2391BF,
32'h3E1378E0,
32'hBE988CB0,
32'h5DF5C8BD,
32'h3EBF27ED,
32'hBEDAB920,
32'h3CDB2844,
32'h3DBBA3E1,
32'hBE283E5F,
32'hBE1A60C3,
32'hBE7B5192,
32'h5DFB3079,
32'h3D2829AA,
32'hBED018BD,
32'h3D60CD11,
32'hBE693315,
32'hBE82C0E4,
32'h3E6FD16C,
32'hBD5B337E,
32'h3E8B8B7A,
32'hBE4FDBA4,
32'hBE08786A,
32'hBD09EB24,
32'h3E60FF0E,
32'hBEA4FD19,
32'h3E05B9B1,
32'h3D800BDE,
32'hBD0CCCAA,
32'hBE8EC626,
32'h3DB61EB6,
32'hBE1CEDD7,
32'hBD71504F,
32'hBE5547AA,
32'hBD33F02E,
32'h3F137830,
32'h3CDF2715,
32'h3ED17111,
32'hBE86CC47,
32'hBE368FBC,
32'hBE8B578E,
32'hBD0EBD71,
32'hBDB1294D,
32'hBD1C2180,
32'hBE0620C4,
32'hBDE0C2D7,
32'h3DF8BC5D,
32'hBE14052C,
32'h3E307BEB,
32'h3E5B4761,
32'hBDF3251C,
32'hBEC4F85A,
32'hBED1118F,
32'hBCFFF5E0,
32'hBDF62F1B,
32'hBE117EAE,
32'h3D84B3B9,
32'hBDA8BFE3,
32'h3DFB16AC,
32'hBDAFC30D,
32'hBE82AEAC,
32'hBEFDE395,
32'h3E209B52,
32'h3D78AF05,
32'h3E385C34,
32'h3EB14D8B,
32'h3DDD1BA0,
32'h3D6FC31B,
32'hBCDB2AE6,
32'hBDAED417,
32'hBC073523,
32'hBE1EFC60,
32'hBD8D06C2,
32'h3D135689,
32'hBDE07496,
32'hBE92DFBB,
32'h3EBEC126,
32'h1DD55F8E,
32'h3E3A041F,
32'h3EA0876E,
32'h3D66A450,
32'hBD77F057,
32'hBE93E43E,
32'hBD59D57C,
32'hBEE4A8F1,
32'hBE14D3B7,
32'hBCE8FCA9,
32'h3D1757F5,
32'hBDA69459,
32'hBDB4363A,
32'hBC134049,
32'hBE91DDA9,
32'hBE65B583,
32'hBE461638,
32'hBE80BAAF,
32'hBE1DFB6B,
32'h3E1798E4,
32'h3DEEAF59,
32'hBE85DBD0,
32'hBD4D1138,
32'h3CD9C308,
32'hBF68E808,
32'h1DC03D7B,
32'h3D8985EC,
32'hBD2D9F80,
32'hBEADC6F0,
32'h3DD5D260,
32'h3E3A148D,
32'h1DC4248A,
32'h3CE0C06E,
32'h3E5E13F3,
32'h3E984E63,
32'h3E27923D,
32'hBDB5DE0A,
32'hBF1D07DD,
32'hBE9B8776,
32'h3D99DEB4,
32'hBEA81F3F,
32'hBE1B878B,
32'h3E9C3FEC,
32'h3DADDB55,
32'hBC9B0640,
32'h3E4E2751,
32'hBEB764C6,
32'hBEA4E139,
32'hBEEF7220,
32'hBCB2ECEE,
32'h3E3B0E9A,
32'hBE3DD3D5,
32'hBE60461E,
32'hBE583671,
32'hBEC8908A,
32'hBD956145,
32'h3D89000B,
32'hBE5963D3,
32'hBE7DB9FE,
32'h3ECDA58A,
32'h3E225455,
32'h3DCE7C2F,
32'hBE0083E9,
32'hBE070FCE,
32'h3DA259A9,
32'h3D538A2D,
32'h3E5F64B2,
32'hBEB0EBD8,
32'hBEAB6AD3,
32'hBE960D4A,
32'hBE37B9A4,
32'hBC4266FD,
32'h3EB116E4,
32'h3D87B492,
32'h3E8DD22F,
32'hBE42C3F1,
32'hBF006870,
32'h3E0989E9,
32'hBD974B03,
32'hBDF10EB4,
32'h3E985C46,
32'hBEA15A58,
32'h3E39DB18,
32'h3E9F39C1,
32'hBEE86774,
32'h3C96313F,
32'hBD59AFB3,
32'hBE510CA8,
32'h3EC35AED,
32'h3EBD074C,
32'hBCA24887,
32'h3E278A5C,
32'h3EC7AAFD,
32'hBCCB9E6B,
32'h3ED02435,
32'h3D8AF17B,
32'h3DA8CED0,
32'hBF4A3D18,
32'hBEC1287B,
32'h3D82F4B1,
32'h3D616257,
32'h3E819BAF,
32'h3EF65CB4,
32'h3EFDAA00,
32'h3EAA12ED,
32'hBE00F18A,
32'hBC9CE299,
32'hBF22D623,
32'h3DA9FB61,
32'h3F0206F9,
32'h3EA352A0,
32'hBF761CD9,
32'h3E14F642,
32'hBF2056F6,
32'hBF87B1B5,
32'h3D41F0AD,
32'hBC6735F0,
32'hBF1C6646,
32'hBD929908,
32'hBE02F247,
32'h3E1A671A,
32'hBEEAEADE,
32'h3EA28D4D,
32'hBF0D4576,
32'h3EA3B6D7,
32'h3EF79CAC,
32'hBE832E41,
32'hBF1998C1,
32'hBEB6B74D,
32'hBEE90DA6,
32'h3EA6756E,
32'h3E55B109,
32'h3EDD39B7,
32'hBF4405A9,
32'h3D5DB680,
32'hBFD00DAA,
32'hBEA1D7D7,
32'hBF1FF081,
32'hBF281C10,
32'h3DF89F7D,
32'h3F0496EF,
32'hC00C4309,
32'h3DF38AB4,
32'hBFB9183A,
32'hBF5B32BD,
32'hBD96FB65,
32'h071E7FA,
32'hBF3831F0,
32'hBE5AFEDE,
32'hBF050B70,
32'hBEE2C020,
32'hBF31EC51,
32'hBECA7D2E,
32'hBF580FDC,
32'hBE5C5913,
32'h3EA460AA,
32'hBC2B02B0,
32'hBF99BB82,
32'hBE58F26D,
32'hBEB54735,
32'h3EB426DD,
32'h3F2C4972,
32'h3E2A811E,
32'hBF624444,
32'hBF4657E3,
32'hC006B8E1,
32'hBF0E280D,
32'hBF85F4ED,
32'hBFF391F2,
32'hBDD9A7E3,
32'h3F072315,
32'hBFAEA710,
32'hBE91B1DF,
32'hBEEB1F7E,
32'hBEB64BA2,
32'h3CDA2AE6,
32'hBD045596,
32'hBEF3BEB8,
32'hBECB245F,
32'hBFB092FA,
32'hBEDB8AA5,
32'hBF8C039F,
32'hBEB468A4,
32'hBF0F84F8,
32'hBE82FE11,
32'hBE5820F9,
32'h3E22A2A8,
32'hBEBB105A,
32'hBDA28244,
32'hBF98484B,
32'hBF8FE876,
32'h3F4C7545,
32'h3D0F195D,
32'hBEF5E265,
32'hBFB2C58E,
32'hBF4E7180,
32'hBF13C9BD,
32'h3E2E6AF8,
32'hBFE14969,
32'h3EBA76FE,
32'h3E5779BC,
32'hBE91FD35,
32'h3EB94F20,
32'h3C1B4F88,
32'h3E481ACB,
32'hBCF51D52,
32'h3D20C0FA,
32'h3EEB3641,
32'h3E10360B,
32'hBEAA3BCC,
32'h3E4E45E6,
32'h3DBB60A2,
32'hBE5E406A,
32'hBEEB9642,
32'h3E93EB33,
32'h3F3B2981,
32'hBE3A425E,
32'hBF099381,
32'hBF00ED03,
32'hBEDF738F,
32'hBEA6E4CA,
32'hBD7335A4,
32'h3F31DE4E,
32'h1DEC7561,
32'hBFA62568,
32'h3E623E60,
32'hBF28A202,
32'h3DD825F2,
32'hBF2E3918,
32'hBF16CF2D,
32'h3F357D98,
32'h3DF48AEB,
32'h3EA71D82,
32'hBDA8CADA,
32'h3E924C97,
32'h3D9B8328,
32'hBD3A09A7,
32'hBEB0EA07,
32'hBD998E30,
32'hBDC2142D,
32'h3EF6269C,
32'h3D4C4D9F,
32'h3E1D50F1,
32'hBE5867DD,
32'hBE9C0A06,
32'hBF391E55,
32'h3F63CA47,
32'hBC494AE1,
32'hBFC56BC6,
32'hBE2AC57A,
32'hBD3E2F86,
32'h3EDF2EC0,
32'h3FBA8E7D,
32'h3DCA7234,
32'hBF4760D8,
32'h3DA68499,
32'h3F0C89BF,
32'h3EA2BEE9,
32'h3E5EAE51,
32'hBCC7DE75,
32'h3D9DE49C,
32'hBC073E81,
32'h3E1CDE1B,
32'h5DE58942,
32'h3D4686A8,
32'h3CB34CE0,
32'hBD44E280,
32'h3EE74353,
32'hBD85A8D2,
32'hBCDAA9B0,
32'hBEE3B33A,
32'h3D48DD03,
32'h3D646514,
32'h3D0D791B,
32'h3E0B3BD7,
32'hBD934B50,
32'h3DC8AF5E,
32'hBDDC2346,
32'h3DA9F0F3,
32'hBE0C24A9,
32'h3DB6F2E7,
32'hBE856D85,
32'h3C6F8045,
32'hBC11660C,
32'h3E421874,
32'hBDDE26AD,
32'h3FB868CE,
32'h3F8F92F7,
32'h3D1A4F07,
32'h3F5E9C80,
32'h3DF21AA0,
32'h3F271E1C,
32'h3F9F3684,
32'h3FBAAB86,
32'hBC83EE40,
32'h3D3198D4,
32'hBC01302E,
32'hBF3323CA,
32'h3EAB5144,
32'h3F369121,
32'hBDE8AC38,
32'h3C963E85,
32'hBE84C4E5,
32'h3F666082,
32'h3E8FDFC0,
32'hBF97CE48,
32'h3EA6F159,
32'hBDE40577,
32'hC004D801,
32'hBEE66266,
32'h4012ECED,
32'hBDA9AA5C,
32'h3F4E331F,
32'hBD44D0F7,
32'hBFDF9094,
32'h3DCE84D1,
32'h3F1AD7FE,
32'hBCFD89AF,
32'h3E76E279,
32'h3E864A60,
32'h3DD8B1CB,
32'hBF63E63E,
32'hBF3CCEC5,
32'hBE81CA8A,
32'h3EF5556F,
32'h3D2E5636,
32'h3DC23EF0,
32'h3E906BFD,
32'hBF96A42D,
32'h3E9F2EEB,
32'hBF324FCF,
32'hBDBD5740,
32'h3E8B95E2,
32'h3F7FB946,
32'h3F097C3D,
32'h3EA0945C,
32'h3C3892DC,
32'h5DD526E3,
32'hBEC8441C,
32'hBDEABE08,
32'h3FD18C4F,
32'hBEF3DC65,
32'hBCC8D1D6,
32'hBE26274C,
32'h3E0CDDE0,
32'h3F8602AE,
32'h3F10D43E,
32'h3F023D68,
32'hBDD4C3ED,
32'h3F4D5261,
32'hBDB0D27B,
32'h3D34F139,
32'h3EADD10B,
32'hBF6F368E,
32'h3EBFC6BA,
32'h3D06719A,
32'h3D21EA54,
32'h3ED9FACE,
32'hBF928AE8,
32'hBDE19B6A,
32'hBE4D69AE,
32'hBF303798,
32'h3F06FA4E,
32'h3E96EF38,
32'h3E299D5F,
32'hBD6AAE75,
32'h3E9B05CC,
32'hBF357BB9,
32'hBED58AE6,
32'h3E0C5FEB,
32'h3F632422,
32'h3E65816A,
32'hBD2069AB,
32'hBE42CD8F,
32'hBF1C1115,
32'h3F2DB75A,
32'hBCA7928D,
32'h3F07AFCC,
32'hBD675477,
32'hBF158AED,
32'hBF2F2342,
32'h3F68AD05,
32'hBE17BA97,
32'hBEEE29FB,
32'hBE1BCA7D,
32'hBDA1FA8E,
32'hBC6C8A29,
32'hBEE921E9,
32'hBE3FB33B,
32'h3E8BAA23,
32'h3E102505,
32'hBD155159,
32'h3F0114B1,
32'hBE918470,
32'h3C6D550F,
32'hBE146550,
32'hBE13E49B,
32'hBF69C869,
32'hBDB74904,
32'h3DFADF3E,
32'h3D3CCF23,
32'h1DDC09D7,
32'h3CC700F0,
32'hBEC6CD85,
32'hBF075D1D,
32'hBDD69BAE,
32'hBC392BAD,
32'hBE4A0612,
32'h3D1F862D,
32'hBF8A8876,
32'hBEA148E1,
32'h3E4FA08C,
32'hBEB642CA,
32'hBF01FE0A,
32'h5DD1A24F,
32'h1DE698E4,
32'hBCAF9ECB,
32'hBE5BD42B,
32'hBDA3D5CA,
32'hBDD45EE0,
32'h3E2F413E,
32'h3DAB3BC1,
32'h3EA9BBB4,
32'hBD72CD48,
32'h3D25AA66,
32'hBDA53181,
32'h3DA3A28F,
32'hBF95CE97,
32'h5DF5B6AB,
32'hBEB83EDA,
32'hBDC2CD88,
32'hBE54C26D,
32'hBF46F42F,
32'h3EB617EB,
32'h3F0A260C,
32'hBEE95FAD,
32'hBE86A129,
32'h3C6BC426,
32'h3E213FBC,
32'hBE844B0E,
32'hBEEB6C50,
32'h3E1B1269,
32'hBDA72791,
32'hBE4A8463,
32'h3CFE6E12,
32'h3D4571D3,
32'h3D403BB7,
32'hBE25F089,
32'hBE6BCE2F,
32'hBE772422,
32'h3E39FBA0,
32'hBF11A2F9,
32'hBCBE7644,
32'h3E43776E,
32'hBDC8EDB2,
32'hBDF6C982,
32'h3D95BFC1,
32'hBFD5F7BB,
32'hBEE4308C,
32'hBE94CCE4,
32'hBE04F769,
32'hBDCE2CB5,
32'hBE06FEDE,
32'h3F18AA23,
32'h3EDC702F,
32'h3E4527D0,
32'hBE6B89B4,
32'h3E817130,
32'hBCF00605,
32'h3C8C4E63,
32'hBE6EAB30,
32'hBDB511F1,
32'hBF1AF541,
32'h3E180CF7,
32'h3D8EC4B6,
32'hBCF89E8C,
32'hBC53334F,
32'h3DB47C2B,
32'h3D92FE9B,
32'h5DE6EF78,
32'h3DAE793A,
32'hBE10E9B5,
32'h3D82800F,
32'h3E7C549E,
32'hBDB13985,
32'h3E6E9A00,
32'hBD93325A,
32'hBE8CDE34,
32'hBE84F56F,
32'h3D7C2024,
32'h3E5867F8,
32'h3E4E091D,
32'h3E0976D6,
32'h3E143DDD,
32'hBC63FD72,
32'h3D917DF6,
32'h3DF721CA,
32'h3DBA830C,
32'h3D63C9AA,
32'h3E875DAE,
32'hBE90C9DB,
32'hBE80C664,
32'hBE1C19EE,
32'hBE00A474,
32'hBF62A346,
32'h3C992D2B,
32'h3C7FD7F8,
32'hBE49879D,
32'hBDE7BC67,
32'h3E4CEEC0,
32'h3DB8B58B,
32'hBD8DE0A8,
32'h3D8F852C,
32'h3E83CD6E,
32'hBDD78F52,
32'h3D4D06A3,
32'h3E12101C,
32'hBC93032B,
32'hBEA97F6E,
32'h3D67098C,
32'h3CFDE655,
32'h1DFB6070,
32'hBE0233BB,
32'h3D5C8BCA,
32'hBF14B24A,
32'h3D057814,
32'hBDA73F70,
32'hBDA9DF48,
32'hBE1B1907,
32'h3D81EDBF,
32'hBE0FA75F,
32'h3D5B335F,
32'hBF46FAD3,
32'hBE2C695D,
32'hBF088A67,
32'hBD379E9F,
32'hBD9F0A0D,
32'hBD97AA5B,
32'h3E28AD48,
32'h3E20B468,
32'hBD073E6F,
32'h3EB33192,
32'h3DF36C21,
32'h3CBAC27E,
32'h3D2621C9,
32'h3E07FABF,
32'h3DFB636D,
32'hBE0382BF,
32'hBDF23B28,
32'h3E610EED,
32'h3E4C5F2F,
32'hBE593291,
32'hBEE2333D,
32'h3C351CE6,
32'hBEF2FB60,
32'hBE406C21,
32'h3E233A25,
32'h3DB0A03C,
32'hBEAC3127,
32'hBE029324,
32'h3D98B0B8,
32'h3EB75AA6,
32'hBF58620D,
32'h3DF64F54,
32'hBE3AB596,
32'hBE2285B1,
32'h3D88E9DF,
32'hBD92998B,
32'h3EEC66F9,
32'hBD4CA613,
32'hBD542C53,
32'h3E5B33C2,
32'h3E05641C,
32'h3DE816A4,
32'hBE2A0188,
32'hBE5CC76B,
32'hBE4D7860,
32'hBF3804B6,
32'hBDD3FC06,
32'h3E835BFB,
32'h3EDDF5D3,
32'hBE22E3BB,
32'hBED1FD3D,
32'h3E383CE6,
32'hBECBC7FF,
32'hBF181F69,
32'hBD1BF010,
32'h3DA71974,
32'hBDB57036,
32'h3D35E6C3,
32'h3EBEF2DE,
32'hBEB56BBC,
32'hBF8F724A,
32'h3DDD118B,
32'hBEAB298C,
32'hBD02D70C,
32'hBCD8468C,
32'hBE942E57,
32'hBE008B5E,
32'hBD27BE67,
32'h3D838905,
32'h3ED9BE26,
32'h3C11FA22,
32'h3E8160B8,
32'hBDFDF89A,
32'hBE43DE74,
32'hBDD13942,
32'hBEE86C05,
32'h3D9B9902,
32'h3EE2662D,
32'h5DE0367F,
32'hBDC1085E,
32'hBE5C278F,
32'h3DB2CE82,
32'hBE95A25A,
32'hBF60657A,
32'h3DA444C8,
32'h3D394914,
32'hBD664FB3,
32'h3C4077B2,
32'h3E7E5C56,
32'hBDDCA914,
32'hBEC91B89,
32'hBDD32691,
32'hBE9C8110,
32'h1DE1DEFB,
32'hBD2F3924,
32'hBE5D64B7,
32'hBE6C4759,
32'hBE66CC0D,
32'hBC6720BE,
32'hBD6BAAA9,
32'h3E722306,
32'h3E475C24,
32'h3E3D0117,
32'hBDCCE18F,
32'h3DBFD420,
32'hBE203BD1,
32'hBDA6E4B1,
32'h3DD81FAD,
32'h3D89FED7,
32'h5CFF4DA,
32'h0EC8E31D,
32'h3D9D86E2,
32'hBE501238,
32'hBF548F8D,
32'hBE5AEEEA,
32'hBDF4AF8F,
32'hBE135908,
32'h3E70B151,
32'h3D267BC2,
32'h3DD2CA56,
32'hBF2A0D1B,
32'h3E265A62,
32'h3E95C0FA,
32'h3C254BEA,
32'h3D962210,
32'hBEA1C81E,
32'hBC630B1B,
32'hBE887D89,
32'hBCA2DC75,
32'hBD87ABDE,
32'hBEA52DF4,
32'hBE0DFC37,
32'h3EA127DD,
32'hBE6C5D78,
32'h3CB95DCA,
32'hBE67D55E,
32'hBD349665,
32'h3DDFC46E,
32'hBE192708,
32'h3E81DE7D,
32'hBE214BEF,
32'h3EEB7455,
32'hBC37254A,
32'hBE7BCE55,
32'hBED88F4F,
32'h3E783267,
32'h3EA72821,
32'h3C99D785,
32'hBE517CA8,
32'hBE107CEA,
32'hBE82C6E9,
32'h3E245BEF,
32'h3F018798,
32'hBD3E69EC,
32'hBCA56D52,
32'hBE6D7811,
32'h3E25A84B,
32'hBE92C471,
32'hBE697763,
32'hBE13F8AE,
32'hBFB307EA,
32'hBD51EB55,
32'hBE531189,
32'h1DC509B1,
32'h3CC13A6E,
32'hBE2BD503,
32'hBEBE0D23,
32'h3E70DFE2,
32'hBDBB9D67,
32'h3DFB75AB,
32'hBEAD07C1,
32'hBE1E669A,
32'hBEF6ED82,
32'h3D9A3205,
32'hBE2CCA26,
32'h3E1E951B,
32'h3EB655F4,
32'hBEB119DF,
32'hBF066541,
32'h3E1783DF,
32'hBCAFF3CC,
32'h3D893029,
32'h3E47B836,
32'hBD33AEDE,
32'hBCB9FCD1,
32'hBE956D25,
32'hBD2A8939,
32'hBE878559,
32'hBD4FB7B4,
32'hBEEE4314,
32'hBF1D7EB9,
32'h3E43E522,
32'hBED3F7F7,
32'h3DEDD090,
32'h3E5B59C9,
32'hBE91053E,
32'hBE564E03,
32'h3E6ED2F2,
32'h3E396D2A,
32'hBCA740C9,
32'hBE2602AD,
32'hBE93E9BC,
32'hBF0389CF,
32'h3E8FC920,
32'h3DBFCC0F,
32'hBD6CDE12,
32'h3F1D6F83,
32'hBE9A16AB,
32'hBE6959CC,
32'h3D9C93C5,
32'hBD7A1BA1,
32'hBE922648,
32'h3D5A55F8,
32'hBDE17771,
32'h3CCDB20B,
32'hBE1B654D,
32'h3D6E2DC0,
32'hBE97958E,
32'hBE42CB10,
32'hBD7CD249,
32'h3E34CEF1,
32'h3CD7AC69,
32'hBF077CD5,
32'hBEB729C7,
32'h3E812028,
32'hBE0D002E,
32'hBCD2FDFA,
32'hBDFEF1B7,
32'h3DA52119,
32'hBDAFC3D4,
32'hBD811CBC,
32'hBE38DB83,
32'hBF030D3F,
32'h3EDCB84B,
32'hBDCB69F3,
32'hBE84F442,
32'h3EF08D01,
32'hBE7834CB,
32'hBE3D880B,
32'h3CF7D6DB,
32'hBD7BE09C,
32'hBEDA2DDF,
32'hBD6876B5,
32'hBDC179A1,
32'hBD9AB753,
32'hBE33AEE0,
32'hBD08FF2E,
32'hBE73784F,
32'hBC93BFBD,
32'h3E9ECFD8,
32'h3EACF3DD,
32'h3E25ADAE,
32'hBE6B97EC,
32'hBE5DBC82,
32'h3E6B2A23,
32'hBD779C9B,
32'h3D3830CF,
32'h3D89289D,
32'h3E0A2349,
32'hBE851A81,
32'hBD72C46B,
32'hBD5E34CC,
32'hBE76588E,
32'hBD909030,
32'h07553B9A,
32'h3CC6AB30,
32'h3EB2D839,
32'h3E780794,
32'h3EE97F1C,
32'hBD30A5A2,
32'h3E24C8D6,
32'hBE64751B,
32'hBE14C0D0,
32'hBD496C45,
32'h3D625B0A,
32'hBE5FCC83,
32'hBCDE3E0E,
32'h3E92E3C5,
32'hBE09EA0E,
32'hBC3E4F8B,
32'h3D98E69F,
32'h3E622F64,
32'hBCB1DDB4,
32'hBE2001E7,
32'hBD84903C,
32'hBF2BB988,
32'hBE22A482,
32'h3DD77E3A,
32'h3ED17F2B,
32'h3D9205B9,
32'hBDC70C69,
32'hBE689C4D,
32'hBEF90F4E,
32'hBD3D2484,
32'hBE84172D,
32'hBD85D729,
32'h3E01F2D6,
32'h3E97F452,
32'h3E9E1D10,
32'h3E278F62,
32'hBCEDA818,
32'h3E70F86F,
32'hBE043F55,
32'h3C35EDA4,
32'h5DE612B8,
32'hBDA1F44C,
32'h3D9D3331,
32'h3E99B302,
32'h3D7C1CA7,
32'h3D079EEB,
32'hBCB6F8F1,
32'hBD40AC1D,
32'hBDE91B4D,
32'hBEACEF91,
32'hBCAC99FC,
32'hBFE0172A,
32'h3C8F39D1,
32'h3E24A1B8,
32'h3E4F6322,
32'h3E3F67AD,
32'h3D78B4D6,
32'hBE40DCBC,
32'hBEF9E799,
32'h3CCF3584,
32'hBF0DACA2,
32'hBE7EC08C,
32'h3E07FDC4,
32'h3DEF8B18,
32'h3F115B12,
32'h3D3120D4,
32'h3DA09CD9,
32'h3D58A29B,
32'hBF87F833,
32'hBDB905BA,
32'hBD82C429,
32'hBE20F352,
32'hBE9F43F7,
32'h3E1BDC3F,
32'h3CB35BE3,
32'hBDE292C0,
32'hBD924295,
32'hBE4AE33D,
32'h3DD6A062,
32'hBE81BE05,
32'h3C582985,
32'hBFE89E27,
32'hBCB2C0B9,
32'hBDC46D3E,
32'hBE04F381,
32'h3E05CADA,
32'h3E27FC9A,
32'hBDAC3B2D,
32'hBDDE1A2B,
32'hBE4ADE7D,
32'h3E45E974,
32'hBE956953,
32'hBE18E3FD,
32'hBDF145D8,
32'h3F1760AE,
32'h3E93676E,
32'h3D333CFA,
32'hBE401C94,
32'hBDF977D3,
32'hBD6D23E2,
32'hBDCFFCEA,
32'h3D974D2F,
32'hBDFA394C,
32'hBCB2D237,
32'h3D522491,
32'h3D8E7711,
32'h3DDB7DBC,
32'h5DFAC04A,
32'h3EBB05D1,
32'hBD89308F,
32'hBD864056,
32'hBF3B6D69,
32'hBD099E80,
32'h3D44C569,
32'h3EA4D397,
32'hBE1D8566,
32'h3A6F778,
32'hBE3976D9,
32'hBCE9A0B7,
32'hBEBFBA3B,
32'hBDFA7069,
32'hBDB50E1E,
32'h3D540254,
32'hBD0A1D09,
32'h3E9BE844,
32'hBE85460B,
32'h3E9CB562,
32'hBCB7129C,
32'hBDADB1AB,
32'hBC3312CD,
32'hBC72CD2B,
32'hBE869127,
32'h3E6AF3B0,
32'h3CC57F57,
32'h3E175300,
32'hBEC5F33F,
32'h3EA64D90,
32'hBE9B025A,
32'hBC9B28B9,
32'h3E16D29C,
32'h3E32AC65,
32'hBE474842,
32'hBE1D452A,
32'h3DBDF7DA,
32'hBE834F6B,
32'h3E9BC751,
32'h3E30842A,
32'hBEB95182,
32'h3E378623,
32'hBE73C926,
32'h3CBAF31B,
32'h3EB8D053,
32'h3EAB9F11,
32'h3DAD7FCA,
32'h3EC09E13,
32'hC02EE412,
32'h5DD2B6DC,
32'hBF2894A4,
32'h3DE9DF6A,
32'h3D305FCD,
32'h3CC4177A,
32'hBEAFA6D1,
32'hBEFF9481,
32'h3E8746CB,
32'hBCCD8483,
32'hBE88BB24,
32'h3E2D1A0B,
32'hBF4E15CF,
32'h3EAD2CD6,
32'h3CD8DE4E,
32'h3E9126EC,
32'hBF4D68E6,
32'hBE0F4A64,
32'hBF0902F9,
32'h3DDC716E,
32'h3F0A6A06,
32'h3E88A804,
32'hBFA03BC5,
32'hBF465007,
32'hBF9C6F94,
32'hBD808F77,
32'hBE95F6E8,
32'hBE93AEB6,
32'hBD9FB71D,
32'h3E91C366,
32'hC03F1BA3,
32'h3EA36E50,
32'hBFCDE5CB,
32'hBF634B3F,
32'h3D99C60B,
32'h3DAE42C6,
32'hBFC1275C,
32'hBF79E1BF,
32'hBFB2B7EC,
32'hBE90F4D3,
32'hBF485FD3,
32'hBF0713AB,
32'hBFAB3BF0,
32'h3EEFF3A2,
32'h3EB742F9,
32'hBC1EAB1F,
32'hBF525909,
32'hBE6B4C5E,
32'hBFA9CA15,
32'h3E6B0E6B,
32'h3F282FA8,
32'h3F3C6D75,
32'hBFA9F312,
32'hBF64BE10,
32'hBFD40AA3,
32'hBEC031AD,
32'hBF62BB21,
32'hBFDCEE8A,
32'h3F2D555B,
32'h3EA5081A,
32'hBFD695C0,
32'h3EAF2BF8,
32'hBF6B39C8,
32'hBF32F882,
32'hBDDD10A6,
32'hBD50BCCB,
32'hBFCD0165,
32'h3E9C980B,
32'hBF488D43,
32'hBEA010A2,
32'hBF9B1574,
32'h3E997DD9,
32'hBFB38D6E,
32'h3E771FEC,
32'h3F03BDC4,
32'h3D6AFD47,
32'hBEF531DB,
32'hBE6C7090,
32'hBF8F2784,
32'hBF51ABB6,
32'h3EAE353F,
32'h3EC7953E,
32'hBE8B29D4,
32'hBF9F9E0F,
32'h3DC3886C,
32'hBF547391,
32'hBE987B14,
32'hBFE3682F,
32'h3EEBEFB6,
32'h3EADB961,
32'hBF0E3C4C,
32'h3DDA82F8,
32'hBDD38D9D,
32'h3EA0ABD6,
32'h3C86E31B,
32'h5DCF518C,
32'hBF1D1B51,
32'hBD21EAD5,
32'hBF42FAC9,
32'h3E11F9CB,
32'h3D54DC4E,
32'hBFC930BE,
32'hBEE18996,
32'hBE64CDE0,
32'hBE8EC988,
32'hBF22A63A,
32'hBE4288EA,
32'hBF26AF69,
32'hBF8A8B13,
32'hBF094E0D,
32'h3E9D6D0F,
32'h3E6EF04B,
32'hBC3102CF,
32'hBF8F0F89,
32'h3E259F76,
32'hBF06D27A,
32'hBE637C8E,
32'hBE99B365,
32'hBD993C4A,
32'h3F22401B,
32'h3E77B71F,
32'hBF3434EC,
32'hBD7B674F,
32'h3DB788BE,
32'h075246AC,
32'h2ED92D5B,
32'hBE2482F5,
32'hBC643CA0,
32'hBDB91A2F,
32'h3F5642A9,
32'h3D44B8B6,
32'hBF6F1B96,
32'hBF20D0D4,
32'hBF67D90D,
32'hBEF143DE,
32'hBF6394BF,
32'hBD92978A,
32'hBEB7CD8E,
32'hBD96A9FD,
32'hBEBED62F,
32'h3CF20EEF,
32'h3E86540C,
32'h3DCDBED6,
32'h3D9DBA61,
32'h3C93DFC5,
32'h3D9744A1,
32'hBD0B8153,
32'h3D6F9911,
32'h3DB380A4,
32'hBD4514B9,
32'h3DCB9EFB,
32'hBC9BDE71,
32'h3D7A157E,
32'h3A18D24,
32'hBCD2A385,
32'hBD793340,
32'h3DBFE82E,
32'hBCE3FBCE,
32'hBC41B02F,
32'hBE2DDC11,
32'h3C036639,
32'hBC88E50D,
32'h3E0E9511,
32'h3DA1C91F,
32'hBDFDE471,
32'hBDA4AB18,
32'h3D4E20E1,
32'hBD7F4417,
32'h0ECBDECB,
32'h3D393D48,
32'hBD7CD204,
32'h3E1988BE,
32'h3C45166D,
32'hBDF0211E,
32'h3D2D64ED,
32'h3FB9AF82,
32'h3EEA2D70,
32'h3D6C3CF7,
32'h3E01A5BC,
32'h3D31469D,
32'h3F4999BE,
32'h3F660B74,
32'hBE8BE8A7,
32'h3D8C919C,
32'h3D7DDFC4,
32'h3DB7FEC8,
32'hBD11C1D8,
32'hBD8A66AD,
32'hBE04FFD2,
32'h3D7994B5,
32'h3D584878,
32'hBE5EA81A,
32'h3F407853,
32'h3E6B7805,
32'hBF9B9625,
32'h3E9ACD0A,
32'hBC2D43FF,
32'hBF9C6A41,
32'hBE5DBB01,
32'h3F7F805E,
32'hBDD4243B,
32'h3F24AE69,
32'h0EC03BCB,
32'hBFC24B5F,
32'h3F110C8A,
32'hBF043D95,
32'h3E87488D,
32'h3EC207C5,
32'h3D3057F9,
32'h1DD35927,
32'hBF0565F2,
32'hBF0AEB62,
32'hBEF8D4AA,
32'h3E35E147,
32'hBDA986A9,
32'h2ECCB7A5,
32'h3EA4B48F,
32'hBF8E457A,
32'h3D847A97,
32'hBF37DD15,
32'hBEA40F84,
32'h3D611B75,
32'h3CAD962D,
32'h3EEADBE2,
32'h3EC6F911,
32'h3F399541,
32'h3D96C01C,
32'h3F06FA54,
32'h3CF2703F,
32'h3DF37DFA,
32'hBE6C72AE,
32'hBC22AF09,
32'hBE990067,
32'h0ED6C75F,
32'h3F42237B,
32'hBD9FD571,
32'hBE95B41B,
32'hBF7E3FCC,
32'h3EE4BBBE,
32'hBEE2DE79,
32'h3F1C7397,
32'h3E968F26,
32'h3EB115B3,
32'hBF17EB9E,
32'h3C0C07C6,
32'h1DF35F38,
32'h3F15486A,
32'hBE672DB9,
32'h3E95922A,
32'hBED73C20,
32'h3F6C9B2B,
32'hBE2DEFF5,
32'h3E75309D,
32'hBE682257,
32'hBF9BE4E4,
32'h3E934AB5,
32'h3E21B866,
32'hBD0B802C,
32'h3F279E4A,
32'h3EC1BE33,
32'h3EDAF4A2,
32'h3D80E532,
32'hBDB0543B,
32'hBFA4E96E,
32'h3EEF0B5B,
32'h3E92CEA4,
32'h3DCEACF2,
32'hBD00D749,
32'hBF5B4EED,
32'hBF4C76FF,
32'h3F349DCF,
32'hBE28CCF2,
32'hBF057F68,
32'hBDBC3BAA,
32'hBD18002C,
32'h3D1E9C0C,
32'hBEFCEE12,
32'h3F132D34,
32'h3E1BA185,
32'hBE45ACBC,
32'h3E596F9A,
32'hBE33AAD2,
32'h3E6C5632,
32'hBED07DA2,
32'hBE388536,
32'hBDE22E63,
32'hBC60E4AF,
32'h3D5D2439,
32'h3E39CE14,
32'h3EA72F3C,
32'hBE553972,
32'h3D9159EB,
32'hBEFD5022,
32'hBF150BC6,
32'h3E7FD64E,
32'h3EBFBA18,
32'h3EC19111,
32'hBE3E15EE,
32'hBE457FA6,
32'hBE01FFAD,
32'h3F22B6B1,
32'hBD9FEC50,
32'h3E347F04,
32'h3E5C46CE,
32'hBD99C16E,
32'hBCE32255,
32'hBEC0738D,
32'hBE5406D7,
32'hBEC6B915,
32'h3E456FA8,
32'hBE5A8AFF,
32'h3ED0D7AD,
32'hBE58B3D7,
32'hBC907AEB,
32'hBF2FD550,
32'hBDDCA024,
32'hBF26AA66,
32'hBD4E3267,
32'hBD3F4FEC,
32'hBDA24E0F,
32'hBDF2C506,
32'hBF42BA32,
32'h3DCD9617,
32'h3E01F1FC,
32'h3F174F2B,
32'h3E86E5AB,
32'h3C16C01F,
32'hBD3074B7,
32'h3C76979E,
32'h3EFAD6DE,
32'h3E5561D0,
32'h3E97B316,
32'hBE709BED,
32'h3EE39335,
32'hBD8BC41A,
32'h5DCA579F,
32'h1DCA13F7,
32'hBF2A82FE,
32'hBCFA28F6,
32'h3E2034B0,
32'hBEEF2B38,
32'hBE36050B,
32'h3ECB4C86,
32'hBE314E6E,
32'hBE9D9CC6,
32'h3EA8D6C1,
32'hBF4D71D1,
32'h3D4CAB9A,
32'h3D294A1B,
32'h3F0AFC2D,
32'h3D96B7AC,
32'hBE485D6A,
32'h3E268322,
32'h3E509442,
32'h3F13FDE7,
32'h3E913483,
32'hBDED453A,
32'hBE8B696A,
32'h3EAE563B,
32'hBEDFB487,
32'hBC1308A5,
32'hBEF84484,
32'h3D57420B,
32'h3E228159,
32'h3C8687B1,
32'hBDDD807A,
32'hBE092578,
32'hBE9D2899,
32'h3DE3E167,
32'h3DEB7377,
32'h3E030BDA,
32'hBDCF00EB,
32'h3E0277A6,
32'hBE72B2CD,
32'h3E0D8D83,
32'h3DDF0EBF,
32'h3DED483A,
32'h3DBDD708,
32'h3E8DAF8D,
32'h3F0C2786,
32'h3D79335D,
32'hBE9BA7DE,
32'hBD3E0635,
32'hBE791ACE,
32'h3EACC2DD,
32'h3D2632D3,
32'hBDCE231B,
32'hBECF9DFB,
32'h3D08658F,
32'hBECBD27E,
32'h3D831B51,
32'hBF41C987,
32'h3DD4161C,
32'h5DC79470,
32'hBC9213C6,
32'h3CEB8FB0,
32'hBD281E50,
32'hBE939549,
32'h3E7D6740,
32'h3E31EBFB,
32'hBDCFBD9A,
32'h3E809C4A,
32'hBE08AFC6,
32'hBCF3217F,
32'h3C5BAEE0,
32'h3ECA714C,
32'h3E8744CA,
32'hBD5D272C,
32'h3E821057,
32'h3D1ACF54,
32'h3D3FF048,
32'hBD32D27A,
32'h3E4BF882,
32'hBDBB172C,
32'h3ECA62F5,
32'h3DFCC12D,
32'h3E81B5F8,
32'hBE13CE66,
32'hBDBFB122,
32'h3E14C397,
32'hBEF63120,
32'hBF67FECD,
32'h3E5C3180,
32'hBE32FB9A,
32'hBDA142F5,
32'hBDB7A827,
32'hBE7FEE10,
32'hBDCF4490,
32'hBEAB0462,
32'h3E03A134,
32'h3D504F3C,
32'h3D903B03,
32'h3CDC959F,
32'h3DC113C2,
32'hBEE2FB2C,
32'h3D1D9C75,
32'hBEA66B1E,
32'hBE205A64,
32'h3E415380,
32'h3ED39D58,
32'h3D494851,
32'hBE168FBB,
32'hBC98C1FD,
32'hBD984665,
32'h3EF35C75,
32'hBE961D39,
32'h3E81D43C,
32'h1DCAC229,
32'hBDA59DB7,
32'hBDB115C5,
32'hBF800A6A,
32'hBF16366C,
32'h3D08F9FB,
32'hBE282B72,
32'hBDFFD976,
32'hBDEF8760,
32'hBE48A973,
32'hBEC2D396,
32'hBEA0CE3C,
32'h3E58BDF9,
32'hBECA2285,
32'hBD1DAE0E,
32'h3D8CF83B,
32'hBE67009E,
32'hBDA71AF6,
32'h3E269C99,
32'h3CEE332B,
32'h3DE8E78A,
32'h3D9113AD,
32'h3E81852B,
32'h3DE1720C,
32'hBE076B50,
32'hBD15890D,
32'hBF1BD4E0,
32'hBECEEF1D,
32'h3D931727,
32'h3E6799A1,
32'hBEA22078,
32'hBDEE5A02,
32'h3E873CF0,
32'hBF4B8308,
32'hBE937DFA,
32'h3E493BF2,
32'hBEC58DD8,
32'h3CECBB14,
32'h41100008,
32'hBEA07DFD,
32'h3E8B3827,
32'hBE2AA6B4,
32'hBD14F55B,
32'hBE9409FE,
32'h3EA3222F,
32'h3C93E768,
32'hBEDFAB14,
32'hBDD0D714,
32'h3D9B01BD,
32'hBF1C6927,
32'hBCB1998B,
32'h3ECFB476,
32'h3E82B76F,
32'h3E13C65E,
32'h3C4D8FD2,
32'h3E66C33D,
32'hBED897A5,
32'hBEF902E4,
32'h3D4F62A6,
32'h3EB5A917,
32'hBDE1EC58,
32'hBDA8B7CB,
32'hBCD4FD9C,
32'hBF3CFB02,
32'hBED34A5F,
32'h3E17E313,
32'hBDBC1EB7,
32'hBD6EBF14,
32'h3CF4592B,
32'hBE1973DD,
32'h3CDB49AE,
32'hBDBC1A04,
32'h3E183F75,
32'hBC8B85A3,
32'h3E90C6A5,
32'h3E8A7105,
32'hBE322815,
32'hBE901D93,
32'h3E8B8B3F,
32'hBDF248DF,
32'h3E25ED89,
32'h3E9D0084,
32'h3EF02441,
32'hBDBC4E51,
32'h3E641436,
32'h3ECC5A81,
32'hBEB22FF5,
32'hBF61CCE9,
32'hBDE0AE7B,
32'h3C9A8069,
32'h3E43F49E,
32'hBE22F505,
32'h3DE7B98F,
32'hBE730341,
32'hBDE6485F,
32'h3E32A5DC,
32'h3EC31DF8,
32'hBD84A599,
32'h3C1D0383,
32'hBDC0F06D,
32'hBEA0B608,
32'hBD93B8D7,
32'hBD2F4E91,
32'hBE174A4B,
32'h3DB21C8E,
32'h5DDF01E9,
32'h3DFEB840,
32'h0ED026CE,
32'h3C1A5FB8,
32'hBDBF4655,
32'h3D8B1DC1,
32'hBE3D5F14,
32'h3EE8B62D,
32'hBE9A89E3,
32'h3E226FD2,
32'h3C87C915,
32'hBE7E018F,
32'hBE93580A,
32'hBD2EE4D9,
32'hBE831A84,
32'h1DC617E9,
32'hBC78DD3C,
32'hBDE988F4,
32'h3C5C1766,
32'hBDFAE22E,
32'h3F09ABF9,
32'h3F329E9D,
32'h3D47E63A,
32'hBDBF2EC0,
32'hBDE1321F,
32'hBE31D439,
32'hBD9808B8,
32'hBDF50580,
32'h5DFB677F,
32'hBFFD134F,
32'h3E6FBF13,
32'hBF29524F,
32'hBE0A8449,
32'h3E5E6432,
32'h3D24C264,
32'hBD8B160F,
32'hBE50B970,
32'h3E4EAC06,
32'hBE2A4A0A,
32'h07543503,
32'hBD9B497D,
32'hBEAB4D45,
32'h3E46465D,
32'hBE3D3DEA,
32'hBE5AC154,
32'h3DA83A3E,
32'hBD845157,
32'hBF3AAD57,
32'h3ECD8496,
32'hBD83EA6E,
32'h3E6A3F69,
32'h3EA7B256,
32'h3D26F983,
32'hBDA5EF48,
32'hBDEF67CF,
32'hBE33C17F,
32'hBE8A7ACF,
32'h5DC4BD5A,
32'h3D700A3E,
32'hBDEF867F,
32'h3E66CF19,
32'hBF03A596,
32'h3E2A845C,
32'h3EEF3C88,
32'hBEBD3F78,
32'hBDA2661D,
32'h3D066012,
32'h3E4462AB,
32'hBE288FE3,
32'h3E7DF715,
32'hBD9524DA,
32'h3E199C79,
32'h3F24DB7A,
32'hBE1CB15B,
32'h3D0F8754,
32'h3DA63134,
32'h3C990E9D,
32'hBF3B5E11,
32'h3E94F7BD,
32'h3DE620E5,
32'hBE040244,
32'h3DC5796A,
32'hBCCAEB59,
32'h3CEF656C,
32'h3E350FCF,
32'h3DC368D0,
32'hBE8C85D6,
32'h3E3ED82B,
32'h3F02B0A0,
32'h3EF97B85,
32'hBD9CF1F0,
32'hBDB37133,
32'hBE108059,
32'h3DF2B743,
32'hBD9A1B22,
32'hBE05ADA2,
32'h3D5DDFB3,
32'h3E0B3E10,
32'hBEB06B2F,
32'h3DFF7347,
32'hBDE06651,
32'hBD8A2EAD,
32'h3DD56D8A,
32'h3DC2758D,
32'h3E5AEEDD,
32'h3DCA3292,
32'h3E3C4641,
32'hBEFE2E88,
32'h3E67256D,
32'hBD92DBBD,
32'hBEB0CD9B,
32'hBEC45FDE,
32'hBD880989,
32'h3D348276,
32'h3D91F9A7,
32'hBD8EAA3B,
32'h3D153434,
32'h3E249134,
32'hBE1BACF0,
32'h3DEC86E0,
32'h3E86D4E9,
32'hBDDC4A95,
32'h0ECA9556,
32'h3E95DC63,
32'hBEF4884C,
32'hBE2BA737,
32'h3E494CF9,
32'h3ED45C0A,
32'hBE7E118B,
32'h3E8BD7A1,
32'hBECA1D50,
32'hBE713A0C,
32'h3DC81A49,
32'h3D4D3139,
32'hBE053E63,
32'h3E8111EE,
32'h3C9CF23E,
32'hBE02C18B,
32'h3E4154CA,
32'h3D044E39,
32'hBE5C7A5E,
32'hBE4BDC15,
32'hBC0AC062,
32'hBD02BFAB,
32'hBE82DD04,
32'h3E4BA039,
32'h3DEB2E45,
32'h3E427879,
32'hBC91738C,
32'hBE007F6A,
32'hBDB0BE30,
32'h3D9B7440,
32'hBE66D9B7,
32'h3D34B0D5,
32'hBFE9B47B,
32'hBE015FD7,
32'h3D74F097,
32'h3E386B40,
32'hBE927873,
32'h3EF16A20,
32'hBDC2994F,
32'hBEC841D0,
32'hBE0656C6,
32'hBDBFDF50,
32'hBEA423C1,
32'h3F17D630,
32'h3E5621E0,
32'h3DD99315,
32'h3E42EBE0,
32'hBDF22DB9,
32'hBE4F1545,
32'hBF04EA5E,
32'hBCF01EA2,
32'h3CCC7A41,
32'hBDC22BF8,
32'h3C989C37,
32'h3F0D315D,
32'h3E0C37CC,
32'hBD4643F7,
32'h3C8A53CA,
32'hBD37E8BA,
32'h3C04B068,
32'h3D9BBDD3,
32'h5DE391C8,
32'hC0044B40,
32'hBC5F861F,
32'hBE221EB3,
32'h3D45EFFE,
32'hBE1EC928,
32'h3DC755EE,
32'h3DC2933E,
32'hBEAA6CAD,
32'hBEC7E5F5,
32'h1DFCEB1F,
32'hBE40BF78,
32'h3EFBCA55,
32'h3E0BB651,
32'h3DEF72E8,
32'h3EB2C7D6,
32'hBD7B08B1,
32'h3E04D248,
32'hBFC280EA,
32'h3CB42AB0,
32'hBCD53F0D,
32'hBD680C57,
32'hBE2DD6FF,
32'h3EA1F879,
32'hBDA465FA,
32'hBF02631E,
32'h3E868840,
32'hBE81AA83,
32'h3EB994A3,
32'h3D3DC1B0,
32'hBE498A50,
32'hBFC42C23,
32'h3D92F9C2,
32'hBCEED657,
32'h3E5F2D1E,
32'hBEC9A418,
32'h1CC942F,
32'hBCB89403,
32'hBE93EB5C,
32'hBDB542A3,
32'h3EC69A70,
32'hBE6FCFEA,
32'h3CA4684F,
32'h3D1588F9,
32'h3EB9B865,
32'hBC58D118,
32'hBD2F5626,
32'hBE1E1791,
32'h3EAA7914,
32'h3CEA0AE8,
32'hBD69388F,
32'hBE7DB265,
32'hBDB3661D,
32'h3EA00C9A,
32'h3E058205,
32'h3D9336BE,
32'h3D742C27,
32'hBE10C799,
32'h3E712D5C,
32'h3E199097,
32'h3D3A4471,
32'hBFB6995B,
32'hBC8E17BC,
32'hBE95B4DB,
32'h3EB64A84,
32'hBEEE7606,
32'h3E298E2C,
32'hBE737A63,
32'hBF0ACF3F,
32'h3E99971C,
32'h3F00B3F7,
32'hBE1BFF9B,
32'h3E203879,
32'h5DCBF12C,
32'h3F13376D,
32'hBD9CBF32,
32'hBD97F72B,
32'hBE5DD72B,
32'hBEDD707F,
32'hBD86FF00,
32'h3CC41077,
32'hBF02E34E,
32'h3D914EBB,
32'hBDD7C68D,
32'h3EA4AA06,
32'h3EDC32B3,
32'h3E1F0126,
32'h3D8E64FD,
32'h3E807025,
32'hBA077F7,
32'h3D7CD34C,
32'hBF51AAAC,
32'hBA52286,
32'h3F248661,
32'h3E1D8A26,
32'h3DAAEC2A,
32'h3F3E2E87,
32'hBEF66F24,
32'hBFAB1EE0,
32'hBEA79A05,
32'h3E821F63,
32'h3E391BBB,
32'h3EE35CE6,
32'hBEA06594,
32'h3E746FCF,
32'hBFD6E092,
32'hBE86D3A9,
32'hBD882041,
32'hBE2F1989,
32'h3C908FA4,
32'h0ED1F7DE,
32'hBE98E3D0,
32'hBE123BDC,
32'h3EFED903,
32'hBDEDDD4B,
32'hBEDBDFA5,
32'hBCB66614,
32'hBE5CA938,
32'h3D29F196,
32'hBD7E109B,
32'hBE26B578,
32'hBF4B4EDF,
32'hBE4DD809,
32'h3EB411D6,
32'h3C04E810,
32'h3EBA09C0,
32'h3F41F7DD,
32'hBF8DF9CA,
32'hBFC121D8,
32'hBFE291D5,
32'h3E4E2CF6,
32'hBF138351,
32'hBE90AB69,
32'h3ED02E0F,
32'h3F2F1C12,
32'hC0431BC0,
32'h3DDF22FB,
32'hBE293983,
32'hBEE2604C,
32'hBDA21590,
32'h3C7CAA71,
32'hBF91C094,
32'hBF872E87,
32'h3E62A929,
32'hBE9303AA,
32'hBEFEE035,
32'hBF6EF75B,
32'hBE883439,
32'h3EBF0CB6,
32'hBD1E201E,
32'hBD5C4BC2,
32'hBE645F25,
32'hBE9BF0C8,
32'hBFF27A7F,
32'hBE7A2F32,
32'h3DF04F90,
32'h3F9561A0,
32'hBFB9797C,
32'hBFBBA55B,
32'hBFB60A9D,
32'h3D9D7DA8,
32'hBF04201F,
32'hC0036EAC,
32'h3E2C32B4,
32'h3ED41B32,
32'hBFC37E1C,
32'hBDD0D051,
32'hBE570972,
32'h3C3F089D,
32'hBD56EDEE,
32'h3CD947A8,
32'hBFC6E4A8,
32'h3EA4DA32,
32'hBF63A7E0,
32'hBE58E791,
32'hBE671886,
32'h3F7E9349,
32'hBF85BAF8,
32'h3EFC8704,
32'hBF59B520,
32'h3F36DF09,
32'hBF365A38,
32'hBE63026A,
32'hBF761041,
32'hBF80D033,
32'h3F8F08E1,
32'h3F3B471A,
32'hBF32EAA5,
32'hC00CDFAC,
32'h3FA50D22,
32'hBF5F24B5,
32'hBE2223F8,
32'hBFD48781,
32'hBFB45531,
32'h3F861C3A,
32'h0ED8A8D8,
32'h3DF905FC,
32'h3EC5A6F7,
32'h3E0B488D,
32'h3D0DF295,
32'h3C89D5C7,
32'hBF3B0010,
32'hBF4E32CC,
32'hBE881AAF,
32'h3EA738DC,
32'hBE8F9A89,
32'hBF0073AA,
32'hBDA8884D,
32'h3DAA48FC,
32'hBF9CDBFE,
32'hBF11BD8D,
32'h3E380A0E,
32'hBE81D729,
32'hBF8470D6,
32'hBE81EC72,
32'h3F4E1C6F,
32'h3C0DE6C6,
32'h3F2D04B7,
32'hBFCCDEA3,
32'h3D9DCA34,
32'hBED190D9,
32'hBE7481C6,
32'h3DBFC002,
32'hBE9AA0EE,
32'h3F75F7BF,
32'hBD691CFB,
32'h3DE506EE,
32'h3EB46026,
32'hBE29D99B,
32'h3C9265DE,
32'h3C4FC230,
32'hBF71C29E,
32'h3D58F5D2,
32'hBDC2F4BB,
32'h3F1BB33C,
32'h3C87B5F8,
32'h3E3934DB,
32'hBE3ABFD5,
32'hBE73701E,
32'hBF30BE27,
32'h3F6B1134,
32'h3D76C62A,
32'hBF7E6857,
32'hBE123A04,
32'hBEB39B1E,
32'h3F8AB666,
32'h3F99A244,
32'h3DD80CC1,
32'hBF8C646A,
32'hBD3B9C72,
32'hBD9BE6A4,
32'hBD664A53,
32'h1DEA1FB9,
32'h3CF16D70,
32'hBDD0911A,
32'hBD1DD7B9,
32'hBD6BA1C6,
32'h3D44E9AE,
32'h3D1AE501,
32'hBD925AED,
32'h3DA3928A,
32'hBCAACB16,
32'h3D250F56,
32'hBDC4E409,
32'hBDD33FED,
32'h3C4551DB,
32'hBCA040B1,
32'h3DB7987C,
32'h3DBF7AC3,
32'hBD88531D,
32'h2E4BB55,
32'hBD683FD2,
32'hBD935650,
32'hBC0B80D3,
32'h3E06EF16,
32'hBE341795,
32'h3DECB06F,
32'h3D043EEC,
32'hBD220BF8,
32'h3F82BBB0,
32'h3F36C665,
32'h3ED19AC5,
32'hBD1F37FD,
32'hBECFD418,
32'hBCD7C6B0,
32'h3E85A43E,
32'hBE7D94CC,
32'hBE31FE33,
32'h3EF6908C,
32'hBC33E3AC,
32'h3D59B4D5,
32'h3D1B4C3D,
32'h3D55ADBF,
32'h3C30EB52,
32'hBE3B9BC6,
32'h3F83A6E4,
32'h3E98BD19,
32'h3F28003A,
32'h3F0941C4,
32'hBEB57262,
32'hBE36B545,
32'h3DBB0EAA,
32'hBF0A9739,
32'hBED7C6FD,
32'h3F03DF72,
32'hBF134AD5,
32'h3E247A4C,
32'h3E5BED22,
32'hBF1FC261,
32'h3DB13551,
32'hBF027B2B,
32'h3CF694EA,
32'h3E5A3D2C,
32'hBD8DCC94,
32'hBDBEE7B8,
32'h3ECB602D,
32'h3E8D0BE7,
32'hBEFDAA0E,
32'h3E1D15E2,
32'hBCE42F7C,
32'hBD5B0FE6,
32'hBE66EF2F,
32'h3E02E8C4,
32'h3D99B744,
32'hBED8C5C3,
32'hBEF8F8C5,
32'hBE8645F9,
32'hBE0BD09A,
32'h3EED0457,
32'hBE9D330E,
32'h3F045901,
32'h3DA952D3,
32'h3F8D4A82,
32'hBF1C5228,
32'hBE04C95C,
32'h3DF28B94,
32'h2EC8CF5D,
32'hBDD7AA4C,
32'hBE02E9A8,
32'h3EB293BB,
32'hBCBAFFE4,
32'hBE36D484,
32'hBFBE25A5,
32'h3E34DE2C,
32'hBED0FE3B,
32'h3F0F2C99,
32'hBD82D81F,
32'h5DF1FC7A,
32'hBF80FC29,
32'hBCF31B99,
32'hBD505E0B,
32'h3E290FE1,
32'h3E18AB90,
32'h3E629B09,
32'hBDA746B0,
32'h3E8CCCD5,
32'h3F10398B,
32'hBDA6D48F,
32'h3E535F77,
32'hBEAB93BF,
32'h3F216CD0,
32'h3E7F0877,
32'h3E33DAB5,
32'h3F4CC0C3,
32'hBF0564B0,
32'h3E769878,
32'h3C0BE39B,
32'hBEB149E8,
32'hBEAEC1D5,
32'h3F7DAF44,
32'h3E2962CF,
32'h3DA53401,
32'hBF05A9D0,
32'hBF263686,
32'hBF220FA7,
32'hBEC707CF,
32'hBE994B86,
32'hBF2736CF,
32'hBE49D829,
32'hBD529790,
32'hBD006B0E,
32'h3DB83331,
32'h3E8895E2,
32'hBD104D58,
32'hBDAD0031,
32'h3F59742C,
32'h3D090918,
32'h3EAA596C,
32'hBECC5305,
32'hBEF0B227,
32'h3EF0C7EB,
32'h3DC8AE24,
32'h3DCFBE5D,
32'h3EBD38E0,
32'h3F275F88,
32'h3E82FAE5,
32'hBEC5DE2B,
32'hBF2366BE,
32'hBED7EC12,
32'h3F1E2045,
32'h3EB60940,
32'h3E54754D,
32'h1DC5D999,
32'h3E688FFE,
32'hBD50412F,
32'hBF86474C,
32'hBD48FA43,
32'h3F89D07A,
32'h3E0BD802,
32'h3DC30098,
32'hBC50D9B5,
32'h3E5AE26A,
32'h3F0A11E1,
32'h3E2480E4,
32'h5DC4DC94,
32'h3EE376FB,
32'h3DC79A1D,
32'h3C6BD2A5,
32'hBD3A6C07,
32'hBF5B3856,
32'hBD964EC4,
32'hBF7BDC3E,
32'hBEF610D8,
32'h3EBFF0E3,
32'h3EC8ED56,
32'h3D1F697F,
32'hBD0FDDF6,
32'h3E38543E,
32'hBEFECE4B,
32'h3ED120FF,
32'h3D9DB0D5,
32'h3C9F4BC1,
32'hBE475A2A,
32'h3E163FA5,
32'hBEEB95B2,
32'hBF3B00F6,
32'h3EAE4ABE,
32'h3E589E4B,
32'hBE4A0DE3,
32'hBDFCCA83,
32'h3DB00058,
32'h3ED67A72,
32'hBF38A1F9,
32'hBEAF5E11,
32'h3E4552E2,
32'hBECF7197,
32'hBF26CEE2,
32'hBE0DFC67,
32'h3DA5F8F1,
32'hBF183F6C,
32'h3EB1FC58,
32'hBF82733D,
32'h3E6AA93D,
32'h3F033603,
32'h3EC57ABA,
32'h3E5C26F5,
32'hBDB19690,
32'hBEB9ACB8,
32'h3D026C47,
32'h3E08CA4B,
32'h3CCD9330,
32'hBE65D1A5,
32'hBE9E02D9,
32'hBE42D39E,
32'h3E3035E0,
32'hBF8B6FB5,
32'hBEAEC4B4,
32'h3E5EAA98,
32'h3DAF324E,
32'hBD2825C3,
32'hBDBDB9F5,
32'hBD10D052,
32'hBF002EAE,
32'h3E2ECD4F,
32'h3E93B311,
32'hBE450D19,
32'h0ECE65AA,
32'h3CC19CCE,
32'hBE91284A,
32'h3D2CB58D,
32'h3E84BDAB,
32'hBE02551F,
32'h3E8ADAAD,
32'h3EBE0BF0,
32'h0757029D,
32'h3D5E2DFD,
32'hBE859EBD,
32'hBF2DD602,
32'hBED3DF21,
32'h3D6B0BEF,
32'hBD86EF23,
32'h3E1A25E4,
32'hBE9A8F1C,
32'hBE0E2F81,
32'hBC99AD8C,
32'hBFFCB9E9,
32'hBEDDAB59,
32'h3DF5128E,
32'hBE8EE935,
32'hBD795BC0,
32'h3D2946F2,
32'hBE9F8BEA,
32'h3E188312,
32'h3E64D36D,
32'h3C560329,
32'hBE71925E,
32'h3D361B85,
32'h3D9B6306,
32'hBD19A294,
32'h3E3B0E83,
32'h3E3FCBF8,
32'hBF0E8880,
32'hBD1CEA84,
32'h3F5984B6,
32'h5CFA6A9,
32'h3D8F8F40,
32'h3E13EAF3,
32'hBF61AAE7,
32'hBEB89B0F,
32'hBE0E3C24,
32'hBC57251D,
32'h3C30DF53,
32'hBDD7A977,
32'hBE020899,
32'h3CFDA349,
32'hBFF1C497,
32'h3E8CA944,
32'h3E99C011,
32'hBEBAF371,
32'hBE00EDE9,
32'hBD9DC44F,
32'hBE67E4B7,
32'h3E643979,
32'hBDBEA461,
32'hBDE214D5,
32'h3D35F5B1,
32'hBD1C2EA6,
32'h3E58F41D,
32'hBE04F01E,
32'hBE42C7EA,
32'h3E2EC4B0,
32'hBE68F11C,
32'h3C10C794,
32'h3EF2F0B8,
32'h3EB30BEE,
32'h3E20BECD,
32'hBDA0745D,
32'hBF2D8775,
32'hBEFE83A7,
32'hBEA342F8,
32'h3CA81B6B,
32'hBD2A5C0D,
32'hBEB8FC65,
32'h3C055F8E,
32'h3CB79E9A,
32'hBF8A232B,
32'h3EB77AC3,
32'h3E6BB948,
32'hBC05C106,
32'hBC5C3FA8,
32'h1DCC9CBA,
32'hBEBE777D,
32'hBE9BE1B3,
32'hBE0FEBCF,
32'h3DF9776D,
32'hBF16B11B,
32'h3C032E6D,
32'hBE12222D,
32'hBD9AF3A5,
32'h3D5E1E6C,
32'h3DA1C18C,
32'hBE84E03C,
32'hBD03340A,
32'h3EDBFCB0,
32'h3E31B7B3,
32'h3CB180CB,
32'h3E4E8D43,
32'hBEAD9CD1,
32'hBF285D83,
32'hBF0C6742,
32'h3F3D4483,
32'hBE076349,
32'hBE8C42F2,
32'hBE28EA42,
32'h3DF73971,
32'hBF289F8C,
32'h3D59FA3C,
32'h3EA039CD,
32'hBE5CD9D4,
32'h2EDA4A48,
32'h3D05205B,
32'hBEB47225,
32'hBEDBC1F4,
32'h3E0FD5BC,
32'hBD532A09,
32'hBF7E0902,
32'h2EC6BAD7,
32'h3DBC1905,
32'hBE124F35,
32'hBE15984E,
32'h3D524E86,
32'hBDA8A41E,
32'hBDF51649,
32'hBE5D36D4,
32'h3E602D9A,
32'hBE3C962B,
32'h3E89C65A,
32'hBEB19851,
32'hBE20A359,
32'hBECF1C64,
32'h3E39D253,
32'hBD67AE38,
32'h3DB68C20,
32'hBE6090CB,
32'hBC2180F3,
32'hBEB487F4,
32'hBDC3041C,
32'h3E143828,
32'hBEE0CF06,
32'hBD9A6E73,
32'h3C4EB1DF,
32'hBF1807E6,
32'hBE097374,
32'h3EC812E6,
32'h3E56AD35,
32'hBE2AC5C3,
32'h3ECCC7C6,
32'h3D66A23F,
32'h3E2FCAB8,
32'hBD377A7C,
32'h3E7CB7FF,
32'hBE811458,
32'h3E7DBF9B,
32'hBF0FC2EB,
32'h3D5AE20C,
32'hBD3A6F7C,
32'h3D875301,
32'hBE871293,
32'hBC8F49D4,
32'hBF3DC61A,
32'h3DCA6B6F,
32'hBEC86D05,
32'hBE8E37ED,
32'hBD914523,
32'h3E99C41B,
32'h3EE7D414,
32'h3E86A98F,
32'hBE1DFF5C,
32'h3F3E517B,
32'hBCF756F1,
32'hBC0A7AA7,
32'hBE8437FD,
32'hBF49E1E4,
32'h3EC506C1,
32'hBE20F532,
32'hBE88FA1C,
32'hBF26303B,
32'hBDC5D2C3,
32'h3DC1AF0C,
32'hBE10F76B,
32'h3E47B5BE,
32'hBE2829D9,
32'h3DAF9F6E,
32'hBFA31146,
32'h3CDA4CDA,
32'hBE9E41EA,
32'h3EA2B2A6,
32'hBF1722EC,
32'hBDB0C23F,
32'hBE1CF331,
32'hBE1DDBE3,
32'hBF5A00AD,
32'h3EC8B47C,
32'hBF2832B2,
32'h1DDB318F,
32'h3F00979F,
32'h3DB6DFA5,
32'h3E49DB3F,
32'h3F1B88AD,
32'hBCFA7662,
32'h3D3BD643,
32'hBD6956BD,
32'hBEEA169C,
32'hBEA6C663,
32'h3E30A352,
32'h3EA4F1AE,
32'hBFF7C1F8,
32'hBD468C10,
32'hBF2365B3,
32'hBE230D27,
32'h3E9B7456,
32'hBEA86771,
32'h3E3147E1,
32'hBF629781,
32'hBEFB064E,
32'hBEAF496A,
32'h3D7A56AE,
32'h3CFE9447,
32'hBDFBEA48,
32'h3EC10FFE,
32'hBDD4AD84,
32'hBED12FB2,
32'h3E8844B3,
32'hBEA0F4F1,
32'hBEAAD13D,
32'h3E5C7EAD,
32'h0EC09FAA,
32'h3E97E121,
32'h3EF1A470,
32'hBE13E5BE,
32'hBDCC6A07,
32'h3D32C947,
32'hBF2C2FF9,
32'hBF24DB9E,
32'h3DD64298,
32'h3D8BCAA6,
32'hBE3ADE14,
32'h3D8EE73B,
32'hBF5A2793,
32'h3E8EB354,
32'h3C9CE46C,
32'hBE97DAB6,
32'h3D233874,
32'hBD972E80,
32'h3DC2307E,
32'hBEF58123,
32'h3E193167,
32'h3E8915B3,
32'h3E0D04BB,
32'h3F17B11E,
32'hBE09B1F9,
32'h5DD585E2,
32'hBD5B6595,
32'hBE46F51B,
32'hBF6E3D5B,
32'h3E10A631,
32'h3D88148E,
32'h3EB62942,
32'h3D2ED93B,
32'hBD2B8CF8,
32'hBDA31057,
32'h3E08D4DF,
32'hBDCE96CE,
32'hBEF5D56B,
32'h3E9D7DB6,
32'h3E7618F7,
32'h3DED92F7,
32'h3EA08E66,
32'hBDD43E79,
32'hBE1FD8A6,
32'hBC00CE53,
32'hBF92CC48,
32'hBD029A98,
32'h1DCE968F,
32'h3E8A8E43,
32'hBEF0E7AF,
32'h3E4D0AE0,
32'h3D8D7F77,
32'h3DB6387F,
32'h3EC0E682,
32'hBE094E25,
32'h3D54F4C2,
32'h3E24CF90,
32'h3E92CEBD,
32'hBF9DCFAD,
32'h5DD1426C,
32'hBDF91225,
32'h3E1FBE18,
32'hBDD4F9C3,
32'h3C596A94,
32'h3CAD302A,
32'h3EEA9BEF,
32'hBDC74173,
32'hBD2A11A0,
32'h3EE4CC55,
32'h3E900EEB,
32'h3E7C2EF6,
32'h3D7AD36E,
32'h3EF398A9,
32'h1DDBACB8,
32'h3C84DB39,
32'hBF9B4DE6,
32'h3E2489E3,
32'hBCE0DF39,
32'h3E94C20E,
32'hBF0596B5,
32'h3E8083EE,
32'h3D8A0741,
32'hBD68042C,
32'h3E27FD73,
32'h3E0F8F39,
32'h3E059280,
32'h3E89EF8F,
32'h3DAE7CE9,
32'hC00C0EFD,
32'h3D41B3D9,
32'hBE8AD238,
32'hBCA38F92,
32'hBEA2230B,
32'h3C098354,
32'hBCA5BDC9,
32'hBD1429CB,
32'h5DCDBCDC,
32'h3E039DAC,
32'h3ED84022,
32'h3DBEE919,
32'hBC1BD7BC,
32'h3CE282A6,
32'h3E6920BB,
32'h3D77DD54,
32'hBDA977FD,
32'hBFC5D1F6,
32'h3D19A44F,
32'h3E15E3EE,
32'h3DEF4E9E,
32'hBE7BEDA0,
32'h3E8F76CC,
32'h3E2B3F6A,
32'hBE890526,
32'hBDDBD597,
32'h3E539A4B,
32'hBE35D447,
32'h3E15713E,
32'h3E93B4E6,
32'hBFD08D1B,
32'h3E292958,
32'h3DFC2BCF,
32'hBE52FD81,
32'hBF92BD13,
32'hBE2E0546,
32'h3C9207A7,
32'hBD7B618C,
32'hBDC7CEBE,
32'h3E02CD72,
32'h3EF1975A,
32'hBD9FAFE2,
32'h3E28990C,
32'hBCEC803A,
32'h3E2A3C6E,
32'hBD0D1BBF,
32'hBD89DB40,
32'hBFB7A48E,
32'hBC606000,
32'h3CC258F0,
32'h3E640B61,
32'hBE9520D2,
32'h3EDB6DD3,
32'h3E7DB5FA,
32'hBEBCBD41,
32'hBEE1E3D8,
32'h3DABF580,
32'hBD9C0968,
32'h3E549E1A,
32'hBC91FD84,
32'hBF1408D5,
32'hBE2308A9,
32'hBD9456DF,
32'hBED985BB,
32'hBF7D0AEC,
32'hBD97213B,
32'h1DC796BF,
32'h3D909A3E,
32'hBE83331D,
32'h3E87ECCF,
32'h3E5C5ECB,
32'hBE580F43,
32'hBE259FDC,
32'hBD50518F,
32'h3E5A3139,
32'h3E037B44,
32'hBE5B091A,
32'hBE5220A6,
32'h3C775032,
32'h3E8A495E,
32'h3E200757,
32'hBEF12864,
32'h3ED3378D,
32'h3E185722,
32'hBEBD43CE,
32'h3ED77CCD,
32'h3E7626C1,
32'hBE98A3FB,
32'h3E9C5403,
32'hBE39B1EF,
32'hBF184CD5,
32'hBEBEDB25,
32'h3E58CBE1,
32'h3D1089FB,
32'hBE855CCE,
32'h075BA6EB,
32'hBCB4B75A,
32'hBD3439E6,
32'hBE014F77,
32'h3EC0A0C7,
32'h3DA217F8,
32'h3E44ECF1,
32'hBE5FD773,
32'hBE84CED5,
32'h3DF77DB5,
32'hBE027D44,
32'hBD756245,
32'hBFBCBCDB,
32'hBD27CCC3,
32'h3E837598,
32'h3D976E8E,
32'hBEA34E48,
32'h3F170653,
32'hBD55E0D1,
32'hBF1D88DD,
32'h3E179663,
32'h3EC3CEBF,
32'hBE549155,
32'h3F0D151E,
32'hBE457468,
32'hBE9015CB,
32'hBE89B51F,
32'h3E542798,
32'h3D5C0855,
32'h3F6BCF26,
32'hBC88EDDA,
32'hBD4D3C17,
32'hBE65C6C2,
32'hBD77BD63,
32'hBE971F7F,
32'h3EE74A30,
32'hBEF37772,
32'hBE33E29B,
32'hBC742A05,
32'hBE63DDF7,
32'hBD512E88,
32'hBE8A8D5E,
32'hBF95C04C,
32'hBE04237D,
32'hBE58F3BD,
32'h3D7A2C62,
32'hBF12E1CB,
32'h3F33E709,
32'hBDCEA2E0,
32'hBF28D67A,
32'hBF4B1009,
32'h3EF64BB1,
32'hBE0E3E70,
32'h3F43EAE5,
32'h3D9A765B,
32'hBF19DE3E,
32'hBFC33885,
32'hBE3AB83D,
32'hBE106199,
32'hBE6D4C67,
32'h3D6856B7,
32'hBC9B3D91,
32'hBED8CF87,
32'hBF696D53,
32'h3E2F135E,
32'h3E8416E3,
32'hBF26EB7E,
32'hBF065364,
32'hBED0021C,
32'hBEE45BCA,
32'hBDD35307,
32'hBDFEF19B,
32'hBF647682,
32'h3E6EECCB,
32'hBF261954,
32'hBEA563E5,
32'h3E313FC8,
32'h3F4CCED6,
32'hBFAD2172,
32'hBFA94ECB,
32'hC0176839,
32'hBE90EC51,
32'h3EEC7A93,
32'hBD802ACC,
32'h3DEE0D16,
32'h3D99F8AD,
32'hBFCC1C87,
32'h3EA24FB9,
32'hBEBFF066,
32'hBF02E128,
32'hBDF40ADC,
32'h1CC3ABB,
32'hBF82B69F,
32'hBF2360C3,
32'h3F47C211,
32'hBEB6B889,
32'hBF10E118,
32'h3F002A46,
32'hBECB6EFF,
32'h3EC916B9,
32'hBF097E87,
32'h3EB25535,
32'hBF020D02,
32'hBE48247F,
32'hBF19AD98,
32'h3E8AF643,
32'h3C9A2FE2,
32'h3F814A74,
32'hBF818368,
32'hBFB19CD3,
32'hBF927D37,
32'h3E9F084B,
32'hBE8D74C3,
32'hBF99ED51,
32'h3E868701,
32'h3E9820E1,
32'hBEF74EB4,
32'h3F126117,
32'hBEB13D2B,
32'h3F216651,
32'hBCF4AF0C,
32'h3D808050,
32'hBF5E34F1,
32'hBE89CEED,
32'hBF078871,
32'hBE12C58C,
32'hBEE2C3F9,
32'h3F525418,
32'h3EDA73BB,
32'h3DA0BFEE,
32'h3ED3F54D,
32'h3EAAA905,
32'hBF4A9D07,
32'hBF126617,
32'h1DC1A279,
32'h3C210B57,
32'hBDA88A1C,
32'h3F799872,
32'hBF2311DF,
32'hBF7DC67A,
32'h3F1BF88E,
32'hBF2A58B6,
32'h3EBDCA59,
32'hBF9FF3AF,
32'hBFB043B1,
32'h3F4C8207,
32'h3E1D75B3,
32'hBEBB9D0E,
32'hBE66651C,
32'hBD9F1EA7,
32'h5DF9D5D4,
32'hBCD82D5C,
32'hBF228C41,
32'h3DB79503,
32'h3EC612F5,
32'hBE48866B,
32'hBE8A3A6A,
32'hBECBC545,
32'hBF543D79,
32'hBDA8446B,
32'hC0031A92,
32'hBDC2BD06,
32'h3E319022,
32'hBEE010E0,
32'h3ECA1F30,
32'hBEE571C3,
32'h3F694E16,
32'h3EE53533,
32'h3EA280ED,
32'hBFA4F1E8,
32'h3F315C20,
32'hBEF033BA,
32'hBE05C178,
32'hBDADC4FD,
32'h3D465A68,
32'h3F8806F7,
32'hBE0B9CF0,
32'h3D144D49,
32'h3DF21675,
32'h3F1851C5,
32'hBD7E4BCC,
32'hBCA3A0F1,
32'hBE5D4642,
32'h3D6D39C0,
32'h5DDA81FD,
32'h3E894071,
32'hBC6BA180,
32'h3E2BD66B,
32'hBE431637,
32'hBDAD9AD2,
32'hBE58208D,
32'h3E0415C6,
32'hBD3AEFE8,
32'hBF191C9D,
32'hBDF5D0AC,
32'hBD4945F5,
32'h3EB05B2A,
32'h3F05F9A4,
32'h3D3601CB,
32'hBEDD837D,
32'h3D4AE9AF,
32'h5DC59E87,
32'h3D25634A,
32'h3DA4C3B5,
32'h3D13BEC5,
32'h2EC9A50D,
32'hBDBCDDEC,
32'hBDA55163,
32'h3D594098,
32'hBC510FEB,
32'hBCA34627,
32'h3DA28DD0,
32'h3D6BCCEF,
32'hBD1B9B93,
32'hBD53A9B1,
32'hBD97A569,
32'hBD3A1CEC,
32'hBCBBBCDA,
32'h3E1CD852,
32'h3E455EAA,
32'hBDA0E3C0,
32'h3CD234EB,
32'hBD32157C,
32'hBDE14537,
32'hBD1F70DE,
32'h3D28D4D9,
32'hBE1A0276,
32'h3E28C3CE,
32'hBD8D1040,
32'hBDBEDF06,
32'h3E27F6FC,
32'h3F433A68,
32'h3E8DE4D9,
32'h3EC4EBDA,
32'hBF16E5F5,
32'hBE1FB886,
32'hBD384C58,
32'h3DC6599E,
32'hBE516C32,
32'h3E5976C2,
32'h1CD1BC9,
32'hBCD196C1,
32'h3F468B59,
32'hBDED2E4E,
32'hBD7554A8,
32'hBF3D3686,
32'h3E58FFCE,
32'hBEB085BC,
32'hBE68B9DA,
32'h3D74CBA1,
32'hBDD0E697,
32'h3F1269AD,
32'hBCCFFC45,
32'h3EBC5E92,
32'hBE6908B2,
32'h3F89D9F9,
32'hBE816F44,
32'h3EAD1297,
32'h3D12CC60,
32'hBE919F02,
32'h3E1C1BD0,
32'h3EF6C1E2,
32'hBE444124,
32'h3DA0C5E1,
32'h3E04FE94,
32'h3E5C84B1,
32'hBED28050,
32'hBD79070E,
32'hBF2A87F4,
32'h3F1A54A5,
32'hBDE7F304,
32'hBD1FC9AB,
32'h3EC3C5F7,
32'hBF0AA30E,
32'hBF16B590,
32'hBD7897DE,
32'hBE90F964,
32'hBED87B57,
32'h3F0E782F,
32'hBEADCF72,
32'hBF295832,
32'h3DD118FD,
32'h3CE98E84,
32'h3F122E52,
32'hBF8AA8D0,
32'h3F0EB97F,
32'hBEECF934,
32'h3EC8AA4D,
32'hBF15918A,
32'hBF066DF6,
32'hBE8C7106,
32'h3F5B95DF,
32'h3DD693D1,
32'hBF854778,
32'hBDE95D4F,
32'h3F3ADEA1,
32'hBF732FCE,
32'h3E90F8E2,
32'h3E89E368,
32'hBF192B19,
32'hBC79FD12,
32'h3CD70E74,
32'hBF6A1B9B,
32'hBECAAF39,
32'h3DC43477,
32'h3EA476D7,
32'h3E7C93DC,
32'h3EE8C9F8,
32'h3F33F75E,
32'hBE6C65E2,
32'hBF7E3315,
32'hBE18EAA9,
32'hBF5D25EB,
32'hBE5B12AD,
32'h3E3946AF,
32'h3E1117BB,
32'h3E1A1243,
32'h3E4143FF,
32'hBF1FABF8,
32'h3E629D47,
32'h3F2D31C7,
32'h3E10F153,
32'h3F146928,
32'hBDCF6DCE,
32'hBED73983,
32'h3F0E5BD7,
32'hBF979BF8,
32'h3E149C6F,
32'hBF573744,
32'hBD5FE356,
32'hBD283D0E,
32'h1CF5C39,
32'hBF18622A,
32'hBEC3F784,
32'h3DC511A3,
32'hBE671FD9,
32'h3F90E5A9,
32'hBDCD42B8,
32'h3E2CB163,
32'hBE208C47,
32'hBEF4B667,
32'h3E375CC3,
32'hBF17314C,
32'h3D667B9E,
32'h3F371F92,
32'h3EE1AA5D,
32'h3F21BE04,
32'hBE83DD4D,
32'hBF5DF682,
32'hBEAEA75C,
32'h2EC04858,
32'h3DFA160B,
32'h3E05F6A1,
32'hBF197EE3,
32'hBE4732DF,
32'hBE0D610B,
32'hBFE689FB,
32'hBE593AE7,
32'h3EE4FE35,
32'h3ECC199E,
32'h3C9CE0C7,
32'h1DE511E3,
32'hBEC32FD4,
32'hBE9A2851,
32'h3DE7A879,
32'h3EADF6F7,
32'h3F374267,
32'h3E54019C,
32'h3E5D25C8,
32'h3D2E8B02,
32'hBE31A297,
32'hBDF6234F,
32'hBEA9D4C8,
32'hBE6AB0A6,
32'h1753A93E,
32'h3DAB8964,
32'hBDE4B481,
32'hBEE9CD6D,
32'hBF46507E,
32'h3DF00DF8,
32'hBE90F8AE,
32'h3C8C5A1E,
32'h3EC8F1F6,
32'hBF0031DD,
32'h3D5FA898,
32'hBCC914EB,
32'hBFC85DE8,
32'hBE7568E5,
32'hBD82FEF4,
32'h3D10843F,
32'hBD82E888,
32'hBDABF5C8,
32'hBDD2E1F8,
32'hBF6CC677,
32'hBE38670D,
32'h3DCEAD04,
32'h3F15F99D,
32'h3D9A8CDD,
32'h3E0D6D01,
32'h3DDA37A9,
32'h3E0A10BF,
32'h3E0ADA62,
32'hBECB356B,
32'h3E7B5B09,
32'h3F393A3E,
32'h3E9245DE,
32'h3E28A4AD,
32'hBE7F9917,
32'hBF6BD1A6,
32'h3D05131B,
32'hBF28F947,
32'h3D0B3C43,
32'h3E90D5C8,
32'h3D3E085E,
32'hBE16371C,
32'h3ED47B14,
32'hBFCF65F9,
32'h3F040305,
32'h3EE16B6C,
32'hBE1100B0,
32'h3CAE69E0,
32'hBD5D545C,
32'hBE514A5C,
32'hBF4B35F3,
32'hBE17A034,
32'h3E51ADCD,
32'h3E826245,
32'h0EC0EC30,
32'h3E8D42C9,
32'h3C96BFE6,
32'hBE1CAC34,
32'hBD68BE75,
32'hBF085D01,
32'hBC4CC3EF,
32'h3F19AC41,
32'hBDA4D6E7,
32'hBC8D70F2,
32'hBDCF4675,
32'hBFAA95A0,
32'h3E1EE4F7,
32'hBF019C99,
32'hBE6A8CF1,
32'h3ED37BC4,
32'hBD410BBD,
32'hBCC62472,
32'h075815E0,
32'hBF9E4EE2,
32'h3F2D5B91,
32'h3EC94A15,
32'hBE974A5D,
32'hBD98BE61,
32'hBD7331A8,
32'hBECFC643,
32'hBFA47F80,
32'hBDE75B8F,
32'h3E849292,
32'hBEAC1719,
32'h0ECED057,
32'h3E6BF739,
32'h3E2AFA49,
32'h3EC1EE8E,
32'hBD906588,
32'hBEB2B5FB,
32'hBE1D29C5,
32'hBDD497F8,
32'hBD866426,
32'hBD699370,
32'h3D758C98,
32'hBFAF3FD6,
32'h3E740CFB,
32'hBDE2E879,
32'h3E750259,
32'h3E331573,
32'hBE8227E3,
32'h3D7F130D,
32'hBEB8C4EA,
32'hBF2A434C,
32'h3E1AF948,
32'h3ED4FF05,
32'hBEC7E0A9,
32'hBC162805,
32'h3CC1DBB9,
32'hBE8E3163,
32'hBFC2BBA8,
32'h3E815CDA,
32'h3DFD7728,
32'hBE083A44,
32'h3E4BEDEE,
32'h3D8E29C6,
32'h1DEB089F,
32'h3E090207,
32'h3D73F53F,
32'h3E6DCA94,
32'hBDB3C4B0,
32'hBFAC8007,
32'h3DBD8715,
32'hBD839483,
32'h3D443846,
32'hBF829185,
32'h5DCAC24D,
32'hBE6E3DBE,
32'h3EC1FB86,
32'h3EB38298,
32'h3D5B9298,
32'h3DF8060C,
32'hBD32C8CC,
32'hBE72A7E6,
32'h3E1D1EE0,
32'h3EE3B93B,
32'hBD5E7A93,
32'h3CE7E025,
32'hBD5DAB2A,
32'h3E7B5387,
32'hBF949F51,
32'h3EFB4404,
32'hBD9D0573,
32'hBEC9F579,
32'h3EAF591B,
32'h3DE39D04,
32'h3E38A238,
32'h3E7F4EA4,
32'hBD9A4E95,
32'h3D39EC7D,
32'hBC39BA44,
32'hC01B3775,
32'h3E38DA52,
32'hBDDBBEE5,
32'h175DD2DA,
32'hBF8F48CA,
32'h3C6715A6,
32'hBEF14417,
32'h3EB28B93,
32'h3EF43BCE,
32'h3DE5F433,
32'h3D8924B4,
32'h3D2D9DBD,
32'h3D9FEF36,
32'h3E6B387C,
32'h3F231634,
32'hBE3E3047,
32'h3D4121BF,
32'h3CF8DA2F,
32'hBE536300,
32'hBF51FDD1,
32'h3EE5CA4E,
32'hBD33A9B9,
32'h3E2996BC,
32'h3DD1CD8D,
32'h3DE2A4B9,
32'h3E20D169,
32'hBE13954D,
32'hBD8F96D1,
32'h3DAC25B6,
32'h3D22A3B6,
32'hC02C04A4,
32'h3EC0B2C9,
32'h3DB2D3DE,
32'hBD7B25F9,
32'hBF3F79CE,
32'hBD48CCF9,
32'h3E0A19C1,
32'h3EF81723,
32'hBF341381,
32'hBEE2D1FD,
32'h3E287281,
32'h3E631B69,
32'h3F0A2059,
32'h3DC166F6,
32'h3EB8D256,
32'hBDDD1EC4,
32'hBDE5DECB,
32'h0EC1302D,
32'hBEEEE530,
32'hBFA40D78,
32'h3EFB1677,
32'hBD28AC4F,
32'hBE1B46C6,
32'h3EA3CBE7,
32'h1DC3746B,
32'h3EC43C7C,
32'h3E5A1D4B,
32'h3E79FD09,
32'h3E614AE0,
32'h3DBCB2D2,
32'hBFE22465,
32'hBDDA27D5,
32'hBD27D51A,
32'h3E23DFCD,
32'hBF2042D0,
32'h3E377AD6,
32'hBEF4D353,
32'h3D1639C0,
32'hBFA46CF8,
32'hBDD5CD02,
32'h3E30AE8B,
32'h3EA8DEB5,
32'h3E9AD78E,
32'h3E916737,
32'h3D9B3738,
32'h3EA0EB0C,
32'hBC485C3F,
32'hBC83D721,
32'hBE0552D7,
32'hBF80F47A,
32'h3C56D486,
32'hBE14A4BC,
32'hBEB076A8,
32'hBF9369CE,
32'hBE10763F,
32'h3E10E68C,
32'hBE884969,
32'h3E144839,
32'hBD51FE24,
32'h3E887764,
32'hBEB4BB91,
32'hBEF45E01,
32'hBD6B277B,
32'h3D4DCC0A,
32'hBECE786D,
32'hBE55AA6D,
32'h3E2D02AB,
32'hBD71A5EC,
32'hBF0855D2,
32'hBEAD4723,
32'hBEFA2E93,
32'hBD9D6A6E,
32'h3EBC5C73,
32'h3EC3E100,
32'h3E779911,
32'h3E9EE83C,
32'h3D06301E,
32'hBDA3F55C,
32'hBE83599C,
32'hBE458D54,
32'hBEBCCFB0,
32'h3E4CE531,
32'hBDDDC0A5,
32'hBF94DEDE,
32'h3E17675F,
32'hBF00F97A,
32'hBE6A68D9,
32'h3D46C962,
32'hBE48B1B3,
32'h3D1045B6,
32'hBE02FC22,
32'h1756BFFD,
32'hBE1768D6,
32'h5DF50904,
32'hBD5F6526,
32'hBDDED7D6,
32'h3F240A23,
32'hBEDCB435,
32'h3E3895D2,
32'hBF34DE8E,
32'hBDF9FE3F,
32'h3E190DB8,
32'h3E0CF6D2,
32'h3F1BD359,
32'hBC3F6EEC,
32'h3EDD7233,
32'hBCEF2C35,
32'hBCEBA427,
32'hBF007F72,
32'hBF172838,
32'hBECAA9BE,
32'h3D31B996,
32'h3E398A6B,
32'hBDEAFDC2,
32'h3EB5ED01,
32'hBF29409B,
32'h3D075C77,
32'hBDA97B03,
32'hBF1111C5,
32'hBE99AE0E,
32'h3E572F0E,
32'h3DE9C025,
32'hBDDB6550,
32'hBEB66B65,
32'hBD85B681,
32'hBDFF423C,
32'h3E64D6AA,
32'hBE532CA9,
32'hBE659B39,
32'hBF7F2394,
32'hBE18584A,
32'hBDC2F782,
32'hBEC06DAE,
32'h3E6F2B0F,
32'h3D5D56A2,
32'h3E660EE6,
32'h2ED4BD29,
32'hBDDFE9BA,
32'h3E170EBF,
32'hBEC5847D,
32'hBF1EB679,
32'h3E8380AB,
32'h3E8E6BC2,
32'h3ECE9C9F,
32'h3D953DF2,
32'h3E800DFF,
32'hBC91AE6A,
32'h3EAEF1BA,
32'hBF4B1687,
32'h3EA3B21C,
32'h3D9C4772,
32'hBD46157B,
32'hBD8E9E1A,
32'hBF040288,
32'h3E352AB3,
32'h3E568481,
32'h3E5C1C8A,
32'h3CD44E24,
32'hBDDDA3A5,
32'hBF6CF3BA,
32'h3E956C3F,
32'hBE31BB1C,
32'hBE053443,
32'h3E222894,
32'h3D011000,
32'hBE8F5ED8,
32'hBD81980E,
32'h3C37D876,
32'h3D71997D,
32'hBEB1764B,
32'hBEB90B1C,
32'h3E365859,
32'h3E16073F,
32'h3DF02D03,
32'h3EAB5B14,
32'h3E5EBD57,
32'hBDBAE302,
32'h3E94D081,
32'hBF246A37,
32'h3D21E71C,
32'h0ED8DEE9,
32'h3EBB4278,
32'hBE8C82B1,
32'hBF0492BA,
32'h3E3DC7DE,
32'hBC4F683D,
32'h3E862F96,
32'h3E8E1E80,
32'hBDF8C3F6,
32'h3E20B78E,
32'h3E6740E6,
32'hBF6850BA,
32'hBCD2D1FB,
32'h3E3B3F3E,
32'h3D302F75,
32'hBED7D6AA,
32'hBD49D833,
32'hBDDC9EEB,
32'hBD7D9454,
32'hBE81B95C,
32'h3E0126B5,
32'h3E87C8B3,
32'h3F00B3E7,
32'h2EC88BE6,
32'h3D4892B2,
32'h3EB3B991,
32'hBE63D290,
32'h3D1B89FD,
32'hBE631C51,
32'hBDCB3747,
32'hBD13E7FA,
32'h3DF05B58,
32'hBDD2B11D,
32'hBF11BDED,
32'h3D918B62,
32'hBE94D798,
32'hBE34311A,
32'h3F10C482,
32'h3E3CAD5D,
32'h3EE7C59B,
32'hBE1758EE,
32'hC0106F97,
32'hBDE4CCC2,
32'h3E841A32,
32'hBE5965FD,
32'hBED953F0,
32'hBD532F1E,
32'h3A1AD46,
32'h3EACF8E4,
32'hBD09C65B,
32'h3E4A0A6F,
32'h3E433841,
32'hBE83B285,
32'hBDD199AB,
32'h3DA7CAF1,
32'h3DD6E3FB,
32'hBE9DE80A,
32'hBE4A5DE2,
32'h3E346C3B,
32'h3E59DDC7,
32'hBE2A0438,
32'h3EA45A89,
32'hBE67C245,
32'hBF069DFF,
32'h3E811917,
32'hBF30253B,
32'h3E73D2E1,
32'h3E214366,
32'h3DADEE5F,
32'h3D90BC58,
32'h3E6371E2,
32'hC00D4A13,
32'hBE63BBC6,
32'h3E5BF337,
32'hBEDDE59D,
32'hBE58DB1E,
32'hBDBE3CB0,
32'hBD89D561,
32'hBE80329C,
32'h3E3242CD,
32'h3CB2A4A7,
32'h3E3812B4,
32'hBE56E1E2,
32'hBE6920A5,
32'h3E0DEE8A,
32'h3DB39BEA,
32'hBE6D5778,
32'hBCA52045,
32'hBEDE2E3A,
32'h3C8135F1,
32'h3EBE32EF,
32'h3EB0907B,
32'hBEF87549,
32'hBE1BCFE0,
32'hBCAF6C68,
32'hBF278CA0,
32'h3D5FBE70,
32'hBDEFF667,
32'hBEC9CA50,
32'h3D967F18,
32'hBCD7F526,
32'hBFDC3BC6,
32'hBF0C6194,
32'h3E3D355D,
32'h3DA5B2B3,
32'h3D9DC6CA,
32'h3D6CE098,
32'h2ED35B6D,
32'h3E4E1385,
32'hBE523D47,
32'h3D3F34E6,
32'h3EE84A41,
32'hBEE739A7,
32'hBE916D95,
32'h3E8050E1,
32'h3E2F0415,
32'h3E95184A,
32'hBD54D490,
32'hBF14F320,
32'h3EB393AB,
32'h3DD3E58A,
32'hBEE42373,
32'hBF0F3FFD,
32'h3E26E031,
32'hBDD1DB46,
32'hBE9669AE,
32'hBF593CE8,
32'h3E06F03C,
32'h3E1F1BD1,
32'h3EC423F3,
32'hBD2DFF18,
32'hBF938E58,
32'hBF90B87A,
32'h3CE6E801,
32'hBE4624D0,
32'h3EB7CA93,
32'hBDDBBFD2,
32'h3D4B0BA7,
32'h3D82DC7A,
32'hBD323305,
32'h3DD777FA,
32'h3F3E38D1,
32'hBFACFF72,
32'hBE4544EB,
32'h3E5F6E5A,
32'hBD42FBCD,
32'h3A1883A,
32'hBE5EDF48,
32'hBF056293,
32'h3E88892A,
32'hBF143210,
32'hBF08D313,
32'hBEDC71B0,
32'h3F5EEAB5,
32'hBE8C7FF0,
32'hBF3D27F0,
32'hBED9F807,
32'h3ECE51D0,
32'h3DEC6156,
32'h3F106813,
32'h3DB83671,
32'hBF29DB23,
32'hBF3E742A,
32'h3DEA6F58,
32'hBF4F91F6,
32'h3F15AA88,
32'h3D897E30,
32'hBCA76121,
32'hBDC7DC52,
32'h3E428755,
32'h3DBE7523,
32'h3E81E556,
32'hBF0E8CD0,
32'hBEFC466B,
32'hBE0EFB8B,
32'hBE0CCC87,
32'hBF4D6BC6,
32'hBD1C1FC5,
32'h3E00CF79,
32'h3E7BA1B1,
32'hBEAB87D7,
32'hBE49C97B,
32'h3DA01CCC,
32'h3FB6DDEB,
32'hBF671B09,
32'hBFA1C610,
32'hBEE8FD3E,
32'hBEA87C02,
32'h3DA5A1EE,
32'h3E47BBDF,
32'hBE50251B,
32'hBE1760E6,
32'h3D90F790,
32'h3DF2EAC5,
32'h3D313569,
32'hBE8A0539,
32'hBCE07B1F,
32'h3D4BA556,
32'hBF66A37C,
32'hBE3CCC6C,
32'hBEF71FA5,
32'h3F29ABA9,
32'hBF0E4D3F,
32'hBF402BC6,
32'hBF4F42C2,
32'hBF9650FC,
32'hBF9960D8,
32'h3ED685DB,
32'hBF1337B5,
32'h3EA647D4,
32'hBEE5437A,
32'hBEEB1E48,
32'h3E69B4EF,
32'h3F7ACF92,
32'hBEFFBD18,
32'hBF9CAB37,
32'h3EAA46FC,
32'hBEED774C,
32'hBDDCF600,
32'hBF6614D0,
32'hBF242E5C,
32'hBF181410,
32'h3EBA77B1,
32'h3F1C5760,
32'h3F6278C6,
32'h3D54997B,
32'h3D6B00BF,
32'hBD0D578B,
32'hBF71D86F,
32'hBE987C53,
32'h3D4CB245,
32'hBE9080AC,
32'h3F381B69,
32'hBE389A28,
32'hBEEB8F25,
32'hBF19090A,
32'hBF61D1E7,
32'h3F485885,
32'hBF446230,
32'hBE9F5FFC,
32'hBF30A5A1,
32'hBEBD7EC6,
32'h3F1B1F0D,
32'h40080C43,
32'h3CA5FD42,
32'hBF3B5520,
32'h3EB00624,
32'hBF2626EE,
32'hBF87D899,
32'hBFC67E55,
32'hBF57DDF1,
32'h3EED3C6B,
32'hBF027C7A,
32'hBFAC1FA0,
32'hBF77AF30,
32'h3EB214ED,
32'h3C87920C,
32'hBCD43348,
32'hBF79D58B,
32'hBFE35724,
32'h3E708F82,
32'h3FB13047,
32'hBEDC9FF0,
32'hBD902C16,
32'hBF950E7C,
32'h3E813FAA,
32'hBFEE8143,
32'hBEDACA80,
32'h3E301EA0,
32'hBF89D9FE,
32'hBF61EBCD,
32'hBF0A1515,
32'h3FA4D293,
32'h3F75AA3F,
32'h3F1066DA,
32'hBF329AFE,
32'h3ED35DA6,
32'hBE6F6CB0,
32'hBE4C6CE9,
32'h3DEF57E7,
32'h3E1857D0,
32'h3F037CCD,
32'hBE95048C,
32'hBCE15033,
32'h3E136E07,
32'h3F89F9D7,
32'h3DD15CA6,
32'hBD99A64D,
32'hBDC1704F,
32'hBDDF60D2,
32'hBD28BF36,
32'hBD7925F1,
32'hBD89534B,
32'hBE044FA6,
32'hBD18874B,
32'h3E599526,
32'h3A1B172,
32'hBE446D91,
32'h1DD9F79C,
32'hBEFF1454,
32'hBEED7EEA,
32'h3C3246D1,
32'hBE48500E,
32'hBE674044,
32'h3CBF9BBC,
32'h3CFB1F49,
32'hBD49E988,
32'hBD8B387A,
32'hBD030428,
32'h3C4C7031,
32'h3CD25207,
32'h3D24D7AE,
32'hBD14C1A7,
32'hBD298294,
32'h3CAAA641,
32'hBD2E5C85,
32'hBD4D75F9,
32'h3D81F511,
32'hBDB7DE04,
32'hBC7720E1,
32'hBC50B544,
32'h3D098302,
32'h3DE4AF0A,
32'h1DFEEE5C,
32'h3CD91447,
32'h3DBC7F15,
32'hBE035BCB,
32'h3D326005,
32'hBD984E69,
32'h2EDD3B11,
32'hBCCD5299,
32'h3C5E4B68,
32'hBDBA10BC,
32'h3D630DE6,
32'hBD931A0F,
32'hBCC47C3E,
32'hBCD821BD,
32'h3EC95571,
32'h3E7CAC3D,
32'h3E5C64D4,
32'h3E595CE9,
32'hBDA870FC,
32'h3C3B8CFA,
32'h3E60148B,
32'hBEADC4F8,
32'h3EA98CBF,
32'hBD31FF54,
32'h3C141644,
32'h3F1BE188,
32'hBF1FFEE2,
32'hBE16CDC9,
32'hBE837E6E,
32'hBDF96650,
32'h3E74BC3E,
32'h3F821943,
32'h3F025E4E,
32'hBD5CBDBB,
32'hBE6906D2,
32'h3DA99F9B,
32'hBF2EF58C,
32'hBF3B0D63,
32'h3F6DD7B3,
32'hBF185352,
32'h3EC2EA2E,
32'hBF23975F,
32'hBEEFE873,
32'hBDC6A5CD,
32'h3DFDCBDD,
32'hBD3283DD,
32'h3D7EB764,
32'h3D93EEC3,
32'h3E8690AB,
32'h3DA3CC99,
32'h3E763C5A,
32'h3E4768DD,
32'h3F1452D1,
32'hBD824FB8,
32'h3CC7F2D2,
32'h3DD2F10E,
32'hBF11E082,
32'hBF423327,
32'h3DE31ED6,
32'hBDF33806,
32'hBE72FBA7,
32'h3E920310,
32'hBE229ED1,
32'hBF026419,
32'hBE54AA47,
32'h3D9949E0,
32'h3E78B5DC,
32'hBF9B9ABB,
32'h3EF5CEDD,
32'hBE9D0860,
32'h3ED3BF16,
32'hBF024488,
32'hBEC4F6DD,
32'h5DE967CA,
32'h3F45732E,
32'h3EC7A604,
32'hBF422F59,
32'hBE4B40FA,
32'h3F01F3A2,
32'hBF84A801,
32'hBD1812E6,
32'h3E347E49,
32'hBF142E52,
32'h3D1C1B6D,
32'h3CC40D59,
32'hBFB1BFCF,
32'hBF71812F,
32'hBF2E1838,
32'h3DA0E310,
32'h3E099010,
32'h3E38621C,
32'h3EDB346D,
32'h3EA55087,
32'hBF3CE91C,
32'hBEDDEADB,
32'hBE7A1395,
32'h3C8FF1D7,
32'hBE202389,
32'h3E47D5E2,
32'hBEEF4B36,
32'h3E1B0E63,
32'hBDF6087A,
32'h3F0668B0,
32'h3E807113,
32'hBD42F6CF,
32'h3F19D820,
32'hBE181845,
32'hBF028B9B,
32'h3DD873F8,
32'hBF372A93,
32'h3D222B14,
32'hBEC8C9A7,
32'hBE2037EE,
32'hBD8D6664,
32'hBD538DC5,
32'hBF2D5E27,
32'hBFD69123,
32'hBF0BDCB4,
32'h3E2945A1,
32'h3F5804BE,
32'hBEBC27D1,
32'h3E832C6A,
32'hBEE40BEF,
32'hBF717654,
32'h3E935728,
32'hBE9B12D4,
32'h3E944169,
32'h3CEF2631,
32'hBEA6060D,
32'h3EA70609,
32'hBF97B721,
32'hBF717988,
32'hBEF9F5D8,
32'hBF14BBCE,
32'h3E09E572,
32'h3ED1C040,
32'hBEEAF531,
32'h3C7F1565,
32'h3E7476E1,
32'hBE810A9F,
32'h3DBAC7EE,
32'h3F008C01,
32'h3ED8D9ED,
32'hBDD967A4,
32'h3CF145BA,
32'hBECC01DD,
32'hBFF65694,
32'hBF3F7241,
32'h3E000A31,
32'h3F364D94,
32'h3E778FB2,
32'h3E81A6C9,
32'hBCAC3AEC,
32'hBF629428,
32'hBDE682A2,
32'hBF05BB52,
32'hBD8C9CAD,
32'h3E562E4D,
32'h3EAC6275,
32'h3D3E4A5F,
32'hBF2284D2,
32'hBFC6E1E6,
32'h3E3B1B0E,
32'hBE220B38,
32'h3E280115,
32'h3E25139E,
32'h3EA8A936,
32'hBDF9B501,
32'hBE33A1F2,
32'hBF619E49,
32'hBE5AB8C9,
32'hBDFF0F9E,
32'hBE86B98B,
32'hBD3F57CC,
32'hBD89827C,
32'hBEA7D16E,
32'hC00AC34A,
32'hBF1DF54D,
32'hBDAF71DF,
32'hBEF0BDD2,
32'h3E4582AA,
32'h3E082059,
32'hBE597A3D,
32'hBE0D774A,
32'hBCC68C68,
32'hBD83018C,
32'h3D8F392F,
32'hBFB4E074,
32'hBF0CD52C,
32'hBD14E893,
32'h3D9A7B0C,
32'hBFC31DE5,
32'h3D401F93,
32'hBF72D036,
32'h3E39DF1E,
32'h3D364043,
32'hBD08D5C6,
32'hBDE63C44,
32'h3EB28ABD,
32'hBF645144,
32'h3ED6C289,
32'hBE0D9B4B,
32'h3D0BB4E8,
32'h3D17270B,
32'h3C6F75DE,
32'hBE66BDC0,
32'hC007445D,
32'hBF7B3E13,
32'h3D9C8C10,
32'hBF5442B5,
32'h0EC68F21,
32'h3D268578,
32'hBDCFEECF,
32'h3D4F7B6D,
32'h3D2C0B0C,
32'hBF0BB725,
32'hBE3362EC,
32'hC00564C9,
32'h3E261AA9,
32'hBDBE2ABB,
32'hBDB629A4,
32'hBF131065,
32'h3D376519,
32'hBF8919E1,
32'h3DBD2220,
32'h3F0B15BF,
32'hBECB2B2A,
32'hBD85027B,
32'hBE2AED44,
32'h3DC4E637,
32'h3EF1F3D8,
32'h3D33EFA1,
32'h3D5C413D,
32'hBCEFB4A4,
32'h3C35DDBC,
32'hBD6BC1B0,
32'hC000D59C,
32'hBCABA31C,
32'h3E04D860,
32'hBF8ABCCC,
32'hBE08EAC9,
32'hBDDC975F,
32'h3E80C6D0,
32'h3E238231,
32'h3E1A3EB9,
32'hBC42D944,
32'h3D7BFE55,
32'hC0608A6F,
32'hBD6DE9ED,
32'hBE164FB5,
32'h3DFD7AAC,
32'hBEF8A761,
32'h3EE5420D,
32'h3D8496B0,
32'h3DAD3D59,
32'h3DCA4DB2,
32'hBD8E9059,
32'hBDB304D2,
32'hBD654666,
32'h3F002917,
32'h3E3B934B,
32'hBDBC5940,
32'h3DD9D415,
32'h3D21FDD5,
32'hBDF1C207,
32'hBE29950E,
32'hC006D973,
32'hBE17CDDF,
32'hBDDFC2B9,
32'h3D1249F3,
32'hBD2CD684,
32'hBDDE037B,
32'h3E89B3FD,
32'h3D2AEAF2,
32'h3E5EE10E,
32'hBE2EA458,
32'h3E293E01,
32'hC044F63E,
32'hBECE4E28,
32'hBCD11E96,
32'h3D88F9E0,
32'hBE69FC0B,
32'h3E4BC489,
32'hBE15B6ED,
32'h3DDF54FE,
32'h3D2A2BBC,
32'h3D8273CA,
32'h3D6D71F3,
32'h3E07388A,
32'h3F2B4FF6,
32'hBCF2F5C6,
32'hBF1F4849,
32'h3D9CC8EB,
32'hBCC4EBD2,
32'hBDD17E31,
32'h3E3D6A1C,
32'hBF73FBDC,
32'hBD3DDC64,
32'hBE425D15,
32'hBE3836FE,
32'h3DFB55E1,
32'hBD7B627F,
32'hBDC95431,
32'h3E791ED9,
32'h3E10F2A5,
32'hBE602AA7,
32'h3C08AC58,
32'hBF8F8E0B,
32'hBE098418,
32'h3DB00BB3,
32'h3E3245F0,
32'hBE9210AB,
32'h3DECEA6D,
32'hBF32D579,
32'h3E8E4032,
32'hBF41930D,
32'h3E954815,
32'hBE0FE022,
32'h3E2FC8F5,
32'h3E75FB10,
32'h1CF771C,
32'hBED15A3E,
32'hBEBA72B5,
32'hBC431811,
32'h3D65391E,
32'hBA0FA85,
32'hBF8EE521,
32'hBEE1B1BC,
32'hBE3C70E7,
32'h3A1BAF1,
32'h3EC403B2,
32'h3E3B05B9,
32'h3DC0EE7B,
32'h3E896F75,
32'hBD66FC99,
32'h3D41F936,
32'h3E27C2EC,
32'h1DC06709,
32'h3E1FF73B,
32'h3D99FAE8,
32'h3D785393,
32'hBD2B4546,
32'h3E56BE2A,
32'hBD4906C7,
32'h3E0FAECB,
32'hC0220D34,
32'hBD0A8F80,
32'hBE658F0E,
32'h3E822208,
32'h3E8C1E7B,
32'h3E0ED90F,
32'hBDFBC9B0,
32'h3D01EBB0,
32'hBC351759,
32'h1DD62A37,
32'hBE86D196,
32'hBF33C752,
32'hBF433447,
32'h3C6299A0,
32'hBF063352,
32'h3EC94A96,
32'hBDF0700A,
32'h3D7EB2EB,
32'h3ED4622E,
32'hBD8DD149,
32'hBD3D7B26,
32'hBC572DD8,
32'h3E5B6B98,
32'hBED7A89F,
32'h3D87AABC,
32'hBE24E891,
32'h3E2D7443,
32'h3EBE3A31,
32'h3D88C0F9,
32'hBF230D78,
32'hBF9FA641,
32'hBE982D57,
32'hBE2BEA8C,
32'h3EA399A6,
32'hBD01B172,
32'h3E87FA83,
32'hBEA4226B,
32'h3E589533,
32'hBE06BAC9,
32'h3CA5B9A0,
32'h3C3D90B9,
32'hBF10CEDB,
32'hBF6F1CAD,
32'h3CC3C5CF,
32'hBEE8D9F9,
32'hBF0B708C,
32'hBF2C3323,
32'hBDB9B50E,
32'h3EAC1C7B,
32'hBDE50B8D,
32'h3E1BBE8A,
32'hBE081275,
32'h3E95653F,
32'hBFC6ABC0,
32'h3E089DF7,
32'hBE172004,
32'h3DED886A,
32'h3E00A732,
32'h3E9FC3A8,
32'hBEBA68BB,
32'hBEB826F7,
32'hBF5D5A6E,
32'hBEC2F747,
32'h3E7B1E91,
32'h3E374DD4,
32'h3E972B22,
32'hBD0EAF4F,
32'h3D4A523A,
32'hBDD6CB9D,
32'h3C96608D,
32'hBD9F1892,
32'hBE84F62C,
32'hBF4264A9,
32'h3E55DA34,
32'hBE976281,
32'hBEF7C456,
32'hBE3348C1,
32'hBF3558AB,
32'h3D82E1E7,
32'h1DC20D33,
32'hBDF0042F,
32'hBE9B463F,
32'h3EA63F7D,
32'hBE57C9F5,
32'h3DB46261,
32'hBF20D1CD,
32'h3D9A1582,
32'hBE81ACE7,
32'h3E573D9C,
32'hBF414BA3,
32'hBE9EA18C,
32'hBF8C588F,
32'h0751471C,
32'h3E80FF26,
32'hBD541201,
32'h3E91A24D,
32'hBE80E2D3,
32'h2EDC66D4,
32'hBD103C39,
32'hBD25BF1B,
32'hBEEA9FE2,
32'hBF4C24A2,
32'hBF135EC5,
32'h3E898C2A,
32'hBD835944,
32'h3CEBED3C,
32'h3F0E2581,
32'hBF42C87B,
32'h3E588FE6,
32'h3EC44060,
32'hBE2F5F1D,
32'hBE4CF2FB,
32'h3E52D86C,
32'h3E432FB1,
32'h3CBBEF96,
32'hBF22A8E7,
32'hBE9A3A7F,
32'hBE1A8497,
32'h3E8AB95B,
32'h3E18C14A,
32'hBCA49229,
32'hBF655B6B,
32'h3E08FD4F,
32'h3DC17893,
32'hBE945D3B,
32'h3E69075C,
32'hBDC717A1,
32'h3E186D3C,
32'hBDCA2561,
32'hBC900331,
32'hBE7CE80E,
32'hBDFEB872,
32'hBEBAC392,
32'h3D1508F3,
32'h3E8965BC,
32'h3DAE97C2,
32'h3E79E753,
32'hBE9CC041,
32'h3E302DC9,
32'hBDA6079A,
32'hBEA5B0D6,
32'hBE32DB2B,
32'h3EAE6CC6,
32'h3DF4317E,
32'h3D8B2538,
32'hBFC65C19,
32'h3D91D26A,
32'hBDCAC83D,
32'h3DEE7D07,
32'hBCDC6CE5,
32'hBD1699D7,
32'hBF3EB775,
32'h3E58BF4A,
32'hBE2F50C8,
32'hBE0D07CA,
32'h3EA2726B,
32'h3C3F69B3,
32'hBE3FEBC7,
32'hBDB1189E,
32'h3D8BDD30,
32'h3E945935,
32'hBE7BF373,
32'hBEC6055E,
32'h3E228F0B,
32'h3E07795C,
32'hBDA4FF62,
32'h3E733AE6,
32'h3E496867,
32'h3D3D3EDB,
32'h3DBB064F,
32'h3E931C21,
32'hBD37261B,
32'hBC6FC9F1,
32'hBEDE5F4E,
32'h3CB877DA,
32'hBFD15935,
32'hBEA05241,
32'h3E079B40,
32'hBE6918AE,
32'h3E1A9F9A,
32'hBE52C5A3,
32'h3D702DF9,
32'h3E37CA31,
32'hBD2AE6E3,
32'hBE1AF724,
32'h3EB0105C,
32'h3E72C347,
32'hBED92619,
32'hBD0EB2EA,
32'h3D84E6FB,
32'hBE2CC102,
32'hBE9C676D,
32'hBEAB5A1F,
32'h3DB0CBD3,
32'h3E2FCE8B,
32'h3E0DEFB3,
32'h3E6D9619,
32'h3E242DB7,
32'hBDC94A13,
32'h3E4A4BFD,
32'h3DEEDBDC,
32'hBE9AEF47,
32'h3E145421,
32'hBE36771A,
32'hBD5911A8,
32'hC003043F,
32'hBDCDE248,
32'h3D0BD898,
32'hBE9866DF,
32'hBE5CE811,
32'h0E5D87A,
32'h3E40B52C,
32'h3DE70956,
32'hBF38D45B,
32'hBF14EF09,
32'hBD971035,
32'hBE3D778D,
32'hBF848C5E,
32'hBE2FBAA9,
32'hBD6FDC17,
32'h3DF90C7E,
32'hBD184999,
32'hBEFB0836,
32'h3E4C89B4,
32'h3DACE2E8,
32'hBD0BB47B,
32'h3C51B12A,
32'h3D883002,
32'hBDC6E536,
32'hBDC1618A,
32'hBF09F18A,
32'hBE16B3B0,
32'hBE589F79,
32'hBDE3686E,
32'hBDEE7C5D,
32'hC015A583,
32'hBEA3BE14,
32'hBEF08F12,
32'hBF10F496,
32'h3DEA6D0A,
32'hBE089D17,
32'hBE0D727D,
32'hBDF2351B,
32'hBF44C6BA,
32'hBDC02EE5,
32'h3E4657FB,
32'h3DFF9DBF,
32'h3E14EC99,
32'hBE01E065,
32'hBC15924B,
32'hBC80793C,
32'h3DC836F2,
32'h3CE45C80,
32'h3E049762,
32'hBEE513E0,
32'hBEA2E397,
32'hBD9A94CE,
32'h3C398E3D,
32'h3CBCC3DC,
32'hBC318712,
32'hBE96EAEF,
32'h3D81E02C,
32'hBDCBE2DA,
32'hBE44DDE8,
32'hBCA73F95,
32'hBFBC785A,
32'hBE9783C4,
32'hBEB9EB37,
32'h3EC645CF,
32'h3E1E8D0C,
32'h1DE25856,
32'h3E75FBEC,
32'h3CBB6E52,
32'hBFA2DAFC,
32'hBE54066C,
32'h3E988695,
32'h3E2A895E,
32'hBD9EAB1E,
32'hBE0E8A14,
32'h3D5C0275,
32'h3E087E9E,
32'h3E062FA2,
32'hBDA24511,
32'h3D542CEC,
32'hBF2031E3,
32'h3DBF5089,
32'h3DB7E2E5,
32'hBD05972F,
32'h3C0E4BD8,
32'hBE451535,
32'hBEABF785,
32'h3C42BEAE,
32'hBE9F56FA,
32'hBEC06CA4,
32'hBDB854E4,
32'hBF69BF55,
32'hBE1DACEF,
32'hBEFBB984,
32'h3DC6112E,
32'hBE0F4AE3,
32'h2ED8C969,
32'h3E54FDFB,
32'h3E94A10E,
32'hBF7A7582,
32'hBF628DA4,
32'hBDE3F273,
32'h3D787F0F,
32'h3EA2480B,
32'hBD269A98,
32'hBD60A08B,
32'h3C68AB2D,
32'h3DB6A737,
32'h3DB35277,
32'h3EDB2769,
32'hBFB2E6FA,
32'h3EA85BE0,
32'h3E9B02AE,
32'hBD3FF45C,
32'hBD80FBC7,
32'hBD88AB44,
32'hBF13B0B4,
32'h3E92DCBB,
32'hBF161F5D,
32'hBE62EF57,
32'hBF024BCF,
32'hBF20A31C,
32'hBE8682E1,
32'hBF2331BC,
32'hBF201CED,
32'hBDCBD605,
32'hBEF8CDE9,
32'h3F015874,
32'hBD02B3D8,
32'hBF2CD452,
32'hBE8071FB,
32'hBEB516AD,
32'hBEA70F6A,
32'h3EE0C839,
32'hBC93264F,
32'h3CA3ACEE,
32'hBD4343DB,
32'hBE563AD8,
32'hBEA5EC73,
32'h3F3BDCC9,
32'hBF40AFB5,
32'hBE4C8151,
32'h3EDC5B13,
32'hBF065D80,
32'h3E017C48,
32'hBE199019,
32'hBE523942,
32'h3EE3C8B3,
32'hBDD45EFE,
32'hBF7E1D85,
32'hBE8DC992,
32'hBF2168B5,
32'hBE9AAB6F,
32'hBECF911E,
32'hBEDC0987,
32'hBE9E8610,
32'hBCE685DB,
32'h3EB815BE,
32'hBFAA7892,
32'h075D31B5,
32'h3F5C5CB3,
32'hBEA88313,
32'h3EF390D5,
32'hBE70E708,
32'h3C40D888,
32'h5DE7D55B,
32'h3E11E0B4,
32'h3E64BF38,
32'hBE58F7E2,
32'h3F102DFC,
32'hBF37C50D,
32'hBDA434C0,
32'hBF6CB5D0,
32'hBF1450E6,
32'h3DA7FAEB,
32'h3E577381,
32'hBF1DE895,
32'h3EB12E4D,
32'h2ECEE9A5,
32'hBF8D91DC,
32'hBEE10AF7,
32'h3F3DE3B2,
32'h3C73E57C,
32'hBE5AE247,
32'hBE6EC10D,
32'hBF1C270A,
32'h3D881F9E,
32'hBEB90A7E,
32'hBE2F47D8,
32'hBEE6806C,
32'h3F9FC169,
32'h3E93C769,
32'h3F7929A6,
32'h3E415952,
32'hBD2F360B,
32'hBCAAF870,
32'hBED78E98,
32'h3E501F4E,
32'h3F062C5F,
32'h3E0247E8,
32'hBEDD8B54,
32'h3F5BD6DB,
32'hBE88EE6D,
32'h3F47735D,
32'h3F18CAB8,
32'h3F0839E0,
32'hBF5166F1,
32'h3D9B1EA3,
32'h3F89B2E3,
32'hBD26B9CB,
32'h3ED9AFCF,
32'h3F770200,
32'h3FC17F7C,
32'h3DC211DD,
32'hBF971C8B,
32'hBEA965BF,
32'h3EF8DDD5,
32'hBF326388,
32'h3EB678D7,
32'hBE03BC01,
32'hBF15680B,
32'h3E98D514,
32'hBCEBAE5A,
32'hBDEEC956,
32'h3CD90F6C,
32'hBCD84E45,
32'hBFC7EBBC,
32'h3EDAAE69,
32'h3FA88909,
32'h3F37BEF1,
32'hBED2E530,
32'hBE294190,
32'hBF480134,
32'h3F0543B6,
32'h1DDFE858,
32'h3F28EE34,
32'hBF9EAD19,
32'hBF49D217,
32'h3E72A947,
32'hBC7ABD23,
32'h3ED0AA45,
32'h3F0A15B6,
32'h3FC73117,
32'hBDE1DCF5,
32'h3C8B5A16,
32'hBDA41B9E,
32'h3D8885C6,
32'h3DAAE1BB,
32'h3D470D55,
32'h3F1777F5,
32'hBE8C6C13,
32'h3E7C64CC,
32'h3F6CAAB5,
32'h3F8AFC56,
32'h3D209636,
32'hBC771F16,
32'h3DC43496,
32'hBE1301E5,
32'h3D008331,
32'h3DB0BC22,
32'hBDCC8C0A,
32'hBEB2CC9E,
32'hBCC3D9D9,
32'h3D0C1DD8,
32'hBE45563A,
32'hBEF36C70,
32'hBDE2D3D0,
32'hBF5C668F,
32'hBF07BA11,
32'h3D36DD8B,
32'hBE780550,
32'h3D3DD175,
32'h3F05B221,
32'hBE879E95,
32'hBDD0B1F5,
32'hBC920122,
32'hBD2893A5,
32'h3C5C5655,
32'hBCB22530,
32'h3D103CBF,
32'h3D1379BC,
32'hBCFFCE25,
32'h3D2EE900,
32'hBE0236BF,
32'h3D5785E0,
32'h3D9C0C99,
32'h1DD08B1C,
32'h3DA30EBB,
32'hBDE727E2,
32'h3DA5F9FA,
32'h3C0A1105,
32'hBDDF1A0E,
32'h3CA44BC8,
32'hBDD50055,
32'hBC0A44AA,
32'hBD65F3C9,
32'hBC2B88F8,
32'hBD32BD93,
32'h3CB0084E,
32'h0ECA2EF8,
32'h3CC21597,
32'hBDBF6262,
32'h3C3E8D6F,
32'h3D123371,
32'h5DED431F,
32'hBD6D9089,
32'hBDDD5C77,
32'h3E3E44CB,
32'hBD6FE74C,
32'hBD151FDB,
32'hBDE4E3CC,
32'h3E7949E5,
32'hBD6FF9ED,
32'h3D08ADC2,
32'hBCCB8456,
32'hBDB694AA,
32'h3F112BAD,
32'hBF084FAE,
32'hBD879031,
32'hBE6B7E4E,
32'hBDEB4061,
32'h3F01494F,
32'h3F17BD66,
32'h3E944C19,
32'h3D34947E,
32'hBE321D87,
32'hBD948E78,
32'hBDFF8C09,
32'hBF0CFBF1,
32'h3E009A67,
32'hBE58D155,
32'h3DA05AD5,
32'hBF0EB74A,
32'hBE51451E,
32'hBEA7E60B,
32'h3F2ED213,
32'h3E5075D8,
32'h3E434832,
32'h3CDA67E0,
32'hBE6D1787,
32'hBF1760CD,
32'h3D4254F9,
32'h3EE86625,
32'h3D65DCA4,
32'hBDA051FF,
32'hBD12986E,
32'hBF5BD4A7,
32'hBEB54753,
32'h3E864FA1,
32'hBC59EC03,
32'h3EB2494A,
32'hBE79DA5C,
32'h3EDA6C1F,
32'hBE2B8C78,
32'hBF647884,
32'h3EBFB61E,
32'hBDEFF15F,
32'hBF15FACB,
32'hBEE5945C,
32'h3F72E8D4,
32'h3E2E850A,
32'h3E8DFE70,
32'hBF0C4CEE,
32'hBF8679F4,
32'h3E32C15D,
32'hBDD237F7,
32'h3F62FFEF,
32'hBF01230A,
32'hBD6F9C6C,
32'hBE2899AA,
32'hBCF1D1DC,
32'h3FADD264,
32'hBF0B11F6,
32'hBE398F30,
32'hBD008421,
32'h3D5A3905,
32'hBFAD08A9,
32'hBF484D24,
32'hBF511C31,
32'hBDC2DD64,
32'h3F297A91,
32'h3CFB33B3,
32'hBD91C2FE,
32'hBF0D146D,
32'hBF43126F,
32'hBE1921EA,
32'hBF04AD29,
32'h3DD49505,
32'hBF80142D,
32'h3C737CFE,
32'hBEDF0BC7,
32'h3D8FF07D,
32'hBE11240C,
32'h3F134FF6,
32'h3E158448,
32'hBEE817B9,
32'hBE4A4458,
32'hBCCCFF0E,
32'hBE6347C6,
32'h3E351786,
32'h3E9529B9,
32'h3F197817,
32'hBE98E94B,
32'h3EBF604E,
32'hBDBE50E0,
32'hBD3EC202,
32'hBE8FA5BC,
32'hBFA5B051,
32'hBF80DBD0,
32'hBD32256A,
32'h3E1820B7,
32'h3D2DCEA6,
32'h3ED054F0,
32'hBE846141,
32'hBF97001D,
32'h3E236D5D,
32'hBEFCA43D,
32'h3F0376E9,
32'hC007257B,
32'hBEA4FE6B,
32'hBF1185B0,
32'hBF943BD2,
32'hBF08B304,
32'hBDC4EAB2,
32'hBFADFFBB,
32'hBD3E4CA1,
32'h3E969C7A,
32'hBDCB52D5,
32'hBEBBD1C3,
32'h3DC59880,
32'hBD913194,
32'h3EF0D628,
32'h3EE54D18,
32'hBEB53461,
32'hBD17B60E,
32'hBDA35FCB,
32'hBE1C7CA7,
32'hBF9876B3,
32'hBF28A357,
32'hBE0108A4,
32'hBEBB7450,
32'h3D98B481,
32'h3E0B84FD,
32'hBCF38028,
32'hBF192DC7,
32'h3D90A02F,
32'hBEF1BDC9,
32'h3E49DF24,
32'hC0117546,
32'h3D83E78B,
32'h3DBF5FB4,
32'h3E293722,
32'hBEAA2C54,
32'h3E657D8C,
32'hBFCF7783,
32'h3C24D581,
32'h3E29A166,
32'h3EC33E3A,
32'hBDA19759,
32'hBD4A12D9,
32'h3E754880,
32'h3D105823,
32'hBEE49915,
32'h3EAF17DD,
32'hBD24A63C,
32'hBD83A092,
32'h3DBC2802,
32'hBF7BEE42,
32'hBFB197CC,
32'hBEF82A10,
32'hBF9556D1,
32'hBDBA362C,
32'h3DB42DFB,
32'hBCB146AF,
32'h3E69510F,
32'hBD115D02,
32'hBE7F00CE,
32'h3C299BA1,
32'hC0189545,
32'hBD58E855,
32'hBE75EDCF,
32'h3ECD5F08,
32'h3F0E65A7,
32'h3E88FEE5,
32'hBEED151F,
32'h3D760719,
32'h3D356C20,
32'h3E876D43,
32'h3DF391EF,
32'h3E6580E9,
32'h3EA97F8B,
32'hBEA9F788,
32'hBF33EFEC,
32'h3F0CE86F,
32'hBDC4F5AF,
32'h3CB50E6B,
32'h3E59BA8F,
32'hBF3E9751,
32'hBFB40CB9,
32'hBE570D68,
32'hBF51114C,
32'hBDA4BE59,
32'h3E3B3D65,
32'h3CA7FF81,
32'hBD363B10,
32'h3D5120CF,
32'hBE7B83EA,
32'h5DFC5517,
32'hC03546A1,
32'h3ECBF06F,
32'hBDBCABBC,
32'h3DE93699,
32'h3EFED9BE,
32'hBEC1E006,
32'hBE9FB689,
32'h3E07E22D,
32'h3DCAD83B,
32'h3DDD0E4D,
32'hBE0E8DED,
32'h3D0E3A60,
32'h3EDB5984,
32'h3C484078,
32'hBF8C3D39,
32'h3CD7CAA7,
32'hBD159780,
32'h3CB25165,
32'h3E22EB1E,
32'hBE7769D5,
32'hBFB4955B,
32'hBE835450,
32'hBF903495,
32'h3E27289E,
32'h3DEB4432,
32'h3E518028,
32'hBD749F14,
32'hBDACA646,
32'hBD44F92B,
32'h3E3B9B3E,
32'hBF822D68,
32'h3F35F1EC,
32'hBD898CD2,
32'h3E49C488,
32'h3E1F2CC3,
32'h3ED49733,
32'hBF4F571A,
32'hBDA19071,
32'h3E315B2C,
32'h3E2336C1,
32'h3D6288B7,
32'h3C9A8AA3,
32'h3EEF3277,
32'h3DC62FFE,
32'hBF46A84C,
32'h3E25F07E,
32'h3C1F4A52,
32'hBCBD6715,
32'hBDE1B062,
32'h3D3744D4,
32'hBF994D23,
32'hBED606D1,
32'hBF2F448D,
32'h3DE51A83,
32'h3C88F983,
32'hBA2A2FD,
32'h3E126E5D,
32'hBE38A20B,
32'hBDD9E3FB,
32'hBDECCA67,
32'hBC59C927,
32'h3DB6BE3A,
32'h3E3DB8CE,
32'h3C620EE6,
32'h3ECC76C3,
32'h3C92F03B,
32'hBF37FB75,
32'h3E47C5C1,
32'hBF7BE0AD,
32'h3EF222D3,
32'hBE8291BD,
32'h3E06BE8B,
32'h3C8440FC,
32'hBD968FE4,
32'hBF546223,
32'hBE507A07,
32'hBD92DE9A,
32'h3D05F905,
32'h3D5C8DB6,
32'hBE694C7F,
32'hBFD37A18,
32'hBE83117E,
32'hBE6BC85D,
32'h3EE30D03,
32'h0EDA76D4,
32'hBD1B2C81,
32'h3EEC6919,
32'hBC05AA08,
32'hBD08E478,
32'hBE2AE26C,
32'h3E2874E5,
32'h3ED911BD,
32'hBE1513E2,
32'h3E94A06C,
32'h3E274590,
32'h3EBEF24D,
32'hBDFB8C62,
32'h3DA0BA4E,
32'hC033B9C2,
32'h3D3B4533,
32'h3D8D2C34,
32'h3E8459AB,
32'hBE1897AB,
32'hBE70555B,
32'hBEB00902,
32'hBEC1D430,
32'hBCC8133C,
32'hBCF9F5FE,
32'h3D5D4DC0,
32'hBDBBEA63,
32'hC0102689,
32'h3E2001D7,
32'hBF0BF907,
32'h3EB734A6,
32'h3DE01D32,
32'h3E678F57,
32'h3E91D40B,
32'h3E4B5B38,
32'hBE2C1125,
32'hBDA53094,
32'h3E312269,
32'h3EF8DAE7,
32'h3E8E0715,
32'h3E7A10C7,
32'h3EAA7D96,
32'h3EC10705,
32'hBECE0194,
32'hBEB1FA64,
32'hBF477336,
32'hBEEDAA18,
32'hBEABB273,
32'h3EA00B78,
32'hBE25D28F,
32'h3D3E25CD,
32'hBEA168AF,
32'hBE286DCC,
32'h3C78C695,
32'h3C9A1524,
32'h1DE96784,
32'h3E0AD1E7,
32'hBFE84BD0,
32'h3E802304,
32'hBE888C40,
32'hBD930F7A,
32'hBE934AF4,
32'h3DE90D5B,
32'h3EC81A03,
32'h3E070EFC,
32'h3E433E0C,
32'hBE80DB55,
32'h3EBD7C4E,
32'hBF357BBD,
32'h3DB9F064,
32'h3E40F7C9,
32'h3EB11392,
32'h3C250201,
32'h3E7DB573,
32'hBF76180B,
32'h3EA3E496,
32'hBF73E037,
32'hBEF2B3BA,
32'h3DF9AD44,
32'h3E2224DF,
32'hBDBCBA6D,
32'hBE0CE9E4,
32'hBEAE9DF5,
32'hBCC0D738,
32'h3D07A61B,
32'h3A76F7C,
32'h3CECF3ED,
32'hBFA2DC0E,
32'h3D892102,
32'h3C5DEA5F,
32'hBEFC71A2,
32'hBE4F57C6,
32'hBE0D4968,
32'h3E033019,
32'h3E0B036D,
32'h3E2BC8A7,
32'hBE5024D6,
32'h3EE0BBCC,
32'hC001546F,
32'hBCCF2146,
32'hBD262641,
32'h3ECB2D1E,
32'hBE6A8E0A,
32'h3E2FCCAE,
32'hBF3654E8,
32'hBE9235DD,
32'hBFB6B8A3,
32'h3CBFF4C0,
32'h3DB0526D,
32'h3EA63ECC,
32'h3E37DC2A,
32'hBD6A2711,
32'h3DC9BB71,
32'hBD8864DD,
32'h3CD20E3D,
32'hBE3F4CD9,
32'hBF1150F6,
32'hBF76B89C,
32'h3E6D971F,
32'hBE06360D,
32'hBE999718,
32'hBD4B2879,
32'hBEC5991B,
32'hBCC6CF72,
32'h3D6FA05A,
32'hBE18E979,
32'hBE2DBA2C,
32'h3D5FF8A6,
32'hBEA06C9D,
32'h3DA87AA5,
32'h3D1A03E8,
32'h3E3645DC,
32'hBEE7F62E,
32'h3E281A1A,
32'hBF1E12C0,
32'hBE00FDAA,
32'hBFA8A4DD,
32'hBC95BD09,
32'h3D886B8A,
32'hBD7C1005,
32'h3E50DDF9,
32'h5DE0D30C,
32'hBDB61734,
32'h3CB150A5,
32'hBCFB7ECC,
32'hBE0830C6,
32'hBF013B4E,
32'hBEC0DC67,
32'h3E806D7E,
32'hBDD49561,
32'hBD62C459,
32'h3E9C473D,
32'hBF451AE1,
32'h3E29723F,
32'h3CDFC016,
32'hBD8471DF,
32'hBE26EBA0,
32'hBE28E7A8,
32'h3DAD1B69,
32'hBE016E7F,
32'hBEACC97A,
32'hBDBA8F8C,
32'hBE308894,
32'h3DC33894,
32'hBDB19F62,
32'hBE1919D4,
32'hBFA7879E,
32'h3E102B92,
32'hBE61F4DF,
32'h3D567FCE,
32'h3E807783,
32'hBEC69257,
32'hBD16AC1B,
32'hBDF5D0CD,
32'h3C3E99F7,
32'hBC64E9B7,
32'hBE2C56C9,
32'hBEDF5D37,
32'h3DA7A2F8,
32'h3D3DF293,
32'hBCB153E6,
32'h3EB3E980,
32'hBE504424,
32'h3E99175A,
32'h3D072943,
32'h3D430BA2,
32'hBD769F0F,
32'h3E113357,
32'h3DEAFEA5,
32'hBDEC47CC,
32'hBEFCD3AB,
32'h3E15C60D,
32'hBD729589,
32'h3D36B2E3,
32'h3DA830EB,
32'h3D131C7F,
32'hBEA9F957,
32'hBCCA7716,
32'hBD4FC3DC,
32'hBC1A4689,
32'hBD5530F1,
32'hBD3590D8,
32'hBEC98FD3,
32'hBD79C08D,
32'h3D0A9E7F,
32'hBC6FCD55,
32'hBEA80C45,
32'hBEB5D95B,
32'h3DDBB96C,
32'h3E78479A,
32'h3D8F05AC,
32'h3ED9E5BE,
32'h3EBAF9ED,
32'h3DA17D25,
32'h3CB5C8D1,
32'h3E34C024,
32'hBE44E26F,
32'h3E2459C2,
32'hBE6CDACC,
32'hBE3CF11C,
32'hBF2BEE22,
32'hBE08B360,
32'h3E94ABD5,
32'hBEDBDA74,
32'hBDAE01BA,
32'hBD4D7C38,
32'hBE1EE525,
32'hBE4E8166,
32'hBD8D6172,
32'hBE2E1440,
32'hBCE72FAB,
32'hBD84C2DB,
32'hBF7552D1,
32'hBE0CD8DD,
32'hBD0C4AA0,
32'hBCF6FE21,
32'hBC758BED,
32'hBEC05EBD,
32'h3DE2C3EC,
32'h3E90AF75,
32'h3D9B3F71,
32'h3E4A0FAC,
32'h3E268A3C,
32'h3CAAB0D7,
32'h3E14C2A7,
32'h3E4D87B0,
32'h3DCF7722,
32'h3D6685C5,
32'hBE7839F9,
32'hBCED93FE,
32'hBFA6A578,
32'hBD7871AE,
32'hBDB46764,
32'hBE880128,
32'hBECB62AD,
32'hBE2DE7F6,
32'hBE7318E1,
32'h3E4B0A56,
32'hBEE5E627,
32'hBF070C75,
32'hBDB84737,
32'h3C68D2E7,
32'hBD141EC7,
32'h3C720B45,
32'hBD8AB896,
32'h3E0AEFEF,
32'h3DA417E2,
32'hBCB41FBE,
32'h3D48D3EC,
32'h3E28E843,
32'h3D0F117C,
32'hBE2499B2,
32'hBE0DA05C,
32'h3D5BD6D1,
32'h3DF0CC6E,
32'h3E130DBE,
32'hBDB8E1BA,
32'hBF0FB7D8,
32'hBF2367B8,
32'h5DF2DA1C,
32'hBFDC396E,
32'hBE9AC5C4,
32'hBE47FFC7,
32'hBEB739AA,
32'hBD7AC2B6,
32'hBE73A96D,
32'hBE899258,
32'h3E470448,
32'hBE4A5EE8,
32'hBE3D27B1,
32'hBE183F58,
32'h3D2516A1,
32'h3E6140FE,
32'h3C04001F,
32'h3D50E6D4,
32'h3C01022D,
32'hBE68A061,
32'hBE7F95C8,
32'h3DC48F72,
32'hBF844629,
32'h3D99FCF2,
32'hBC95D39E,
32'hBE44351A,
32'h3F26E969,
32'h3E57D941,
32'hBCC9D777,
32'hBD588AC5,
32'hBEBE544E,
32'hBEBF2C2C,
32'h3DC5AD36,
32'hC006B338,
32'hBE5F6A02,
32'hBE3DAC82,
32'h3F24881E,
32'h3E5028F7,
32'hBD18AE3C,
32'h3DD2F499,
32'h3D1D5A14,
32'hBE4B745F,
32'hBE05EE5F,
32'hBE47BD73,
32'hBF12A7CB,
32'hBE6D2A79,
32'h3D28DC61,
32'hBC56B029,
32'h3E967A3F,
32'hBE62EA11,
32'hBDC9354B,
32'h3E06144F,
32'hBFB46D2B,
32'h3EF7B39F,
32'h3EBDDE8D,
32'h3D64F702,
32'h3DD1D21B,
32'h3E9C659D,
32'h3E770D12,
32'hBDA489A2,
32'h3EB7FDAC,
32'h3D7BDB71,
32'h3D8726E7,
32'hC037A401,
32'h3D847BFF,
32'hBE7DD029,
32'h3E645E67,
32'hBECA1AA2,
32'hBECC0240,
32'h3E05A5B1,
32'h3E6B478A,
32'hBF00149C,
32'hBEEE90C4,
32'hBEB8DB2F,
32'hBF00941D,
32'hBF3DDEA1,
32'hBD7DF89C,
32'hBD08AA9D,
32'h3E66DBDF,
32'hBCC66A54,
32'h3D1CF724,
32'h3E51595F,
32'hBFAB1D62,
32'h3D5B305A,
32'h3C1571CF,
32'hBECC6472,
32'hBE453921,
32'h3EA05075,
32'h3D80C31F,
32'h3F1FFB9F,
32'hBCAA4ADA,
32'hBF183943,
32'hBF0E41A0,
32'hC01B3C80,
32'hBCF6BE1E,
32'hBD55D867,
32'h3E39AF21,
32'hBF11FCD6,
32'hBE79775B,
32'h3EEB7F7C,
32'hBE71540B,
32'hBF13BAC5,
32'hBE52FD8B,
32'hBF23952A,
32'h3DABB962,
32'hBF834D3B,
32'h2ED04F75,
32'hBDC0B377,
32'h3F1F3016,
32'hBE090400,
32'hBE06B9AB,
32'h3ECFC59B,
32'hBF47F1F0,
32'hBE2FF95A,
32'hBF3067F6,
32'hBF5FDBC6,
32'h2ECE70E2,
32'h3D778671,
32'hBF408360,
32'h3F357BE4,
32'h3E5C3D8F,
32'hBF2A431C,
32'hBEDA3EE6,
32'hC004CFE6,
32'h3EE66E54,
32'h0EC7BFBF,
32'h3EE789BB,
32'hBE43161B,
32'h3DDD1D9A,
32'h3EC4B17D,
32'hBEDD0D73,
32'hBE7051B9,
32'h3E9E4C5F,
32'hBF5312F9,
32'h3E3823BE,
32'hBF5C4B6F,
32'h3D3870A7,
32'hBC109891,
32'h3F1AC12F,
32'h3F1723E0,
32'h3F0573E5,
32'h3EADB698,
32'hBF6E1782,
32'h3E90596A,
32'hBF46D169,
32'hBE61292C,
32'h3EF73DBD,
32'h3C74B09B,
32'hBF73B01B,
32'h3ED74850,
32'h3DAA3597,
32'hBF0B1C92,
32'hBF1C6554,
32'hBF5CAAA7,
32'h3ECAE15A,
32'h3DADD7EE,
32'h3F2BEEE6,
32'h3E355220,
32'h3F2EB887,
32'hBEB25D3D,
32'h3F1457D9,
32'hBED69D11,
32'h3F1642D6,
32'hBF05FC3E,
32'h3F5B6BE3,
32'hBF1B744D,
32'hBD7BABB8,
32'h3DEC3473,
32'h3DD16193,
32'h3F963607,
32'h3F111836,
32'h3F2D7BC6,
32'hBF2916AF,
32'h3EC14603,
32'hBF576028,
32'h3EE12246,
32'h3EDD2C55,
32'hBED8BCEF,
32'hBF852421,
32'h3EA7C356,
32'h3ECC70E5,
32'h3E6BE6B1,
32'hBDB9DFCD,
32'h3C214F82,
32'h3F820997,
32'hBE0BCC3D,
32'hBF7C71D4,
32'hBE98D168,
32'h3F19AAB2,
32'hBF2936A5,
32'h3F1880DE,
32'hBE94F7B1,
32'h3DF5FCB1,
32'h3E52094E,
32'h3F2BAB48,
32'h3E364748,
32'hBC90A06F,
32'h3DC71FF3,
32'hBE6EA9E6,
32'h3F0D8A25,
32'h3DBF9BED,
32'h3EEA7E98,
32'h3E8D9B7C,
32'h175C31B3,
32'hBEE390B0,
32'h3DCFDAE1,
32'h3EDD6C2B,
32'hBDA15326,
32'hBF9136C3,
32'hBDBC1A8E,
32'h3F1A3AA9,
32'hBE0A623E,
32'h3E3D2A4D,
32'hBD3E525A,
32'h3FB1C951,
32'h3D750FE0,
32'h3D8A83B7,
32'h3D0A85B3,
32'h3EE17303,
32'h3E29A302,
32'h3D854660,
32'hBE0E2592,
32'h3D1EF216,
32'h3EA2E8DD,
32'h3ED32555,
32'h3D78B491,
32'hBCA2598E,
32'hBDA2BDF4,
32'h3E1B26AC,
32'h3E959E6E,
32'h3D5FED48,
32'hBE9CAB7C,
32'h3E90F510,
32'h2EDC9CCD,
32'hBE3C895B,
32'hBD6CE51B,
32'hBE481D91,
32'hBD059B84,
32'hBDA9F02E,
32'h3D418A1E,
32'hBDE89270,
32'h3D2C3EF0,
32'h3DF6CBDE,
32'h3D2E5D2C,
32'h3F2D21CC,
32'hBE0505DB,
32'h3DA67D27,
32'hBC506D34,
32'h3CD90F07,
32'hBD39DB6F,
32'hBDCA27DB,
32'h3F28CFD3,
32'h3E847F8E,
32'hBCCE338B,
32'h3D8F528B,
32'h075A64A6,
32'hBC236FE4,
32'h3D04AF12,
32'hBD8DA0AC,
32'hBD6FE039,
32'hBCCDD64B,
32'hBEA5C4E6,
32'h3D7123A2,
32'h17542812,
32'hBDB1A705,
32'hBDA7EA8F,
32'h3D861720,
32'h3F059487,
32'hBD73D899,
32'h3D40F91D,
32'hBD2C8CA1,
32'hBDC9986B,
32'h3F743B68,
32'hBCBACE79,
32'hBDA6191E,
32'h3CBD58EB,
32'h3C9DB0C3,
32'h3E139F17,
32'hBC2C276E,
32'hBD876F4B,
32'h3D60682E,
32'h3D13E01D,
32'h3F0A40EE,
32'h3E270C83,
32'hBDAC523E,
32'h5DD72113,
32'h3CB744C3,
32'h3DB8411F,
32'hBE1980DD,
32'hBECAE663,
32'hBD49BF35,
32'hBEBBFD91,
32'hBD9F3B1F,
32'hBD28B6CF,
32'h3E9634B2,
32'h3E1FC115,
32'hBD0830A6,
32'h3E0590B7,
32'hBD0313FC,
32'hBE47D3F7,
32'h3F00FA50,
32'h3E1E428D,
32'hBDEC4AC3,
32'h3DF7D96C,
32'hBD469DDF,
32'hBC19BF59,
32'h3EC2FCA6,
32'h3F9566EA,
32'h3D97194E,
32'h3E0C872E,
32'hBD06F72F,
32'hBD74BAF0,
32'hBE83E120,
32'h3F2C08FF,
32'hBE4608B5,
32'hBD2F8AF3,
32'h3CA5DF91,
32'hBDD3F6FF,
32'h3EC6A34A,
32'hBF59A595,
32'hBDD6FF92,
32'hBEEED04C,
32'h3F1D93F1,
32'hBED04548,
32'hBE4EF1F0,
32'hBE0E2613,
32'hBE64DD32,
32'h3F469612,
32'h3D8609AC,
32'hBEB48FE6,
32'hBF10FFDC,
32'h3F21CEDE,
32'h3EF08CAE,
32'h3F2E0532,
32'hBF059210,
32'hBF2FC3D2,
32'h3EA03F54,
32'h3EBC2027,
32'h3F0A4318,
32'hBF253AE9,
32'hBD9AB5EB,
32'h3D1AE89D,
32'h3E432C5B,
32'h3F43E370,
32'hBF67E2CA,
32'hBE413DDA,
32'h3CCF1E9B,
32'h3D3B7EBE,
32'hBF82FE7A,
32'hBDD2DDBA,
32'hBF1FFBF3,
32'h3F1E01B5,
32'h3F08F543,
32'h3E7D9165,
32'h3E1E5424,
32'hBF1C1635,
32'hBF8ABD17,
32'hBF082E3A,
32'hBE922C68,
32'hBE5C6A51,
32'hBF93DAC5,
32'h3F119488,
32'h3DFBF100,
32'hBCAE2BF3,
32'h3F0F9465,
32'h3DC766E1,
32'hBDF0F4ED,
32'hBEBD2ABC,
32'hBEEC9F28,
32'hBEE1E727,
32'h3D26D78F,
32'hBE59B166,
32'hBD2C98F0,
32'h3F2744FC,
32'hBF931CD0,
32'h3F65ABE0,
32'hBD9878E9,
32'hBD48A803,
32'hBE25393F,
32'h3E74A071,
32'hBEA8AD0A,
32'h3EF152D6,
32'hBE891748,
32'hBE294A72,
32'h3EEF85D9,
32'hBE85E6F5,
32'hBF42EF58,
32'h3EA492AE,
32'hBE61D913,
32'h3EA1AC46,
32'hBFCD77BC,
32'hBE9FEB35,
32'hBE54B45A,
32'hBD463CC3,
32'hBE32CDFB,
32'h3F065A2D,
32'hBF163095,
32'hBCE8201D,
32'hBF23C78E,
32'h3E4F14C3,
32'h3C36B63C,
32'hBEABFF6C,
32'hBE94DF77,
32'h3EE260DA,
32'hBF81DCAD,
32'h3DD64EF9,
32'hBC8F6B45,
32'h3D2E3AC9,
32'h3E6BBE7C,
32'hBF3DEA12,
32'hBF7F61B4,
32'hBE86C02D,
32'hBFA13F0A,
32'h3F35A6F9,
32'h3E34F87F,
32'h3E51C791,
32'hBD22E8A2,
32'h3DAA0B9B,
32'h3E835D4E,
32'h3CE80E5B,
32'hBF8014DE,
32'h3EF0767F,
32'hBEEF6A45,
32'h3EDB432D,
32'h3EDFFEF8,
32'h3F0A464B,
32'hBEC19CD9,
32'hBD26E914,
32'h3F036251,
32'h3F07D583,
32'h3DF3B252,
32'hBE961BDF,
32'h3E64AFF6,
32'hBEBDF0EF,
32'hC001C2B5,
32'hBE8FED27,
32'h5DCB03DA,
32'hBDC92A56,
32'h3E5D84AA,
32'h3E932692,
32'hBFA12B2B,
32'hBEB34238,
32'hBFCB9576,
32'h3DB59C6D,
32'hBE70BDF3,
32'hBE240FA8,
32'h5DF8392C,
32'h3EB788F5,
32'h3E4F331F,
32'h3E97D4CC,
32'hBFA654BF,
32'h3CCC4CB4,
32'hBE445B7B,
32'h3E0FB77B,
32'h3F501E66,
32'h3EB26A42,
32'h3EEC2AC8,
32'hBE9CAD6C,
32'hBDC2ECD6,
32'h3EDC4F10,
32'h3E9582D7,
32'hBE3D4AFC,
32'h3DF0E484,
32'hBF047BFF,
32'hBF993CBD,
32'hBD2861EA,
32'hBC5CF3C3,
32'h17585695,
32'h3E020395,
32'h3EFCA280,
32'hBF8F8F93,
32'hBE21FFF8,
32'hBF6763E2,
32'h3EC0E172,
32'h3D67A414,
32'h3D979E57,
32'h3E90E9E2,
32'h3DE655E3,
32'h3F014C94,
32'h3E954D26,
32'hBE3CE3F5,
32'h3E3C632F,
32'hBDF54709,
32'hBC746AAF,
32'h3F3F582E,
32'h3E5D816E,
32'h3E5E3610,
32'h5DF86305,
32'hBFC068FA,
32'h3ECDA888,
32'hBDAB5EEC,
32'hBE20CFFB,
32'hBC50321E,
32'hBDC8E900,
32'hBF8F1FD8,
32'h3F4A86B0,
32'hBC42ACF6,
32'h3C82AFC9,
32'h3E9FAD5F,
32'h3EBC6A9B,
32'hBFD15A45,
32'hBDCB90C3,
32'hBEBB01CF,
32'h3E162595,
32'hBE117198,
32'h3D2900FA,
32'h3E530200,
32'h3E5308F9,
32'h3F221C8C,
32'h3E5CE9DD,
32'h3E481725,
32'h0ED24596,
32'hBD875B35,
32'h3D344903,
32'h3E838D5A,
32'h3E94C882,
32'hBED2074F,
32'h3E2282CD,
32'hC002A502,
32'h3E1B1678,
32'h3E181490,
32'hBDD72588,
32'hBE9B0599,
32'hBC18A816,
32'hBF4F6F45,
32'h3DE02CDB,
32'hBCD50DEA,
32'hBD5D6B93,
32'h3DDA301C,
32'h3F407F77,
32'hBFB92686,
32'hBD307194,
32'hBF566F79,
32'h3EC5BE18,
32'hBD7095B5,
32'h3E867B65,
32'h3E54E2B1,
32'h3E938406,
32'h3DCC74A5,
32'h3DE1CDE7,
32'h3E3C07E3,
32'h3D33F496,
32'hBEA18018,
32'h3DEC30EB,
32'h3E780B28,
32'h3ED228F0,
32'hBEC29FD2,
32'h3DD5BBC1,
32'hC0068344,
32'h3E26D593,
32'hBEA91EED,
32'h3E5C7108,
32'hBE84A0BF,
32'hBD88B7B0,
32'hBD38F2B6,
32'hBF6716D9,
32'hBD95D2DA,
32'hBDB595B4,
32'hBD2DB3E4,
32'h3DC18CD5,
32'hBFC0C46D,
32'h175CF894,
32'hBE7DC786,
32'h3E9217F2,
32'h3DD3A204,
32'h3D30F1D5,
32'hBD2574DE,
32'h3E136C52,
32'h3E16E054,
32'h3DD8A013,
32'h3DCA8B62,
32'hBE9D0D12,
32'hBD7261FE,
32'h3E1F495D,
32'h3EC6B2CA,
32'h3ED30CB5,
32'h3CE243EB,
32'h3E9A1E3E,
32'hBEFA129D,
32'h3DEC2988,
32'hBE4714CF,
32'hBDEBE607,
32'hBE7AD9F2,
32'h5DF21CE1,
32'hBD0213F0,
32'hBEB51B8D,
32'hBCA48B83,
32'h3CC2D4C1,
32'h3D465519,
32'h3E79FB16,
32'hBED4C869,
32'h3DAA3201,
32'hBE0F295C,
32'h3E466D5E,
32'h3D8758B9,
32'h3DB34548,
32'h3EA16E0B,
32'h5DF21C28,
32'hBDC6D310,
32'h3E13D64A,
32'h3EA098A5,
32'hBF206993,
32'h3E11E45B,
32'h3E193584,
32'h3EE0D4DA,
32'h3F249B64,
32'hBE3C8C3F,
32'hBE7452AB,
32'hBE1231DE,
32'hBECFEFC3,
32'hBEA86549,
32'h3D8B3E7C,
32'hBD925E67,
32'h3DB0844B,
32'hBDCEA37E,
32'hBE85C312,
32'h3D9D38F4,
32'hBD8FAC71,
32'h3E43E4D6,
32'h3ED51AC3,
32'hBE864BB8,
32'h3E2FB269,
32'hBE762038,
32'hBE0B4E64,
32'hBE46DD48,
32'hBD8FCCA5,
32'h3E5DDF39,
32'hBCBBAA37,
32'h3EC9A09E,
32'h3E48493C,
32'h3E4F616D,
32'hBF4C3B5C,
32'h3DE74FB9,
32'h3CAEA131,
32'h3E2D912C,
32'h3DAEAF78,
32'h3E08D471,
32'hC001E785,
32'hBE1C73C1,
32'hBF481FB2,
32'hBDE9AB15,
32'h3D9437D9,
32'hBD93DE12,
32'h3D9FA151,
32'hBD87E46B,
32'hBE9209FF,
32'hBD0B2CD0,
32'h5DCBA710,
32'h3E2A28D3,
32'h3E416AC1,
32'hBF5F5FDB,
32'h3E855EFF,
32'h3D154091,
32'hBE2A4870,
32'h3D9B4571,
32'hBEBF0AB6,
32'h3D7381B8,
32'h3D5CAF82,
32'hBDC56E0D,
32'h3D2777B7,
32'h3E3A2320,
32'hBFC53488,
32'hBD9295F3,
32'hBD2D9B2A,
32'h3DE83C5F,
32'hBE9D4CF0,
32'h3E686EBA,
32'hBF80DED4,
32'hBE3E2641,
32'hBF86E237,
32'h3E432F4B,
32'h3E3BA373,
32'h3EB2469D,
32'h3CAB5197,
32'hBE55F90C,
32'h3EA23191,
32'hBD59EFF9,
32'hBCD109FC,
32'hBD6BD420,
32'h3E3986CD,
32'hBF558469,
32'h3E871016,
32'h3DC98C0E,
32'h3DBBE1EB,
32'h3DD0762C,
32'hBF083860,
32'hBD4CE650,
32'h3CFE22A3,
32'hBEA69E78,
32'hBE07B458,
32'h3EEAA802,
32'hBE75AD66,
32'hBD73FB35,
32'hBE8CE354,
32'hBD4D7A8A,
32'hBF173566,
32'hBD67AAE7,
32'hBED8E64D,
32'hBE73A86C,
32'hBF810AA9,
32'h3EB33301,
32'h3D244CE9,
32'h3E8B28FF,
32'hBC0578D2,
32'hBE42C5E9,
32'hBD18D881,
32'hBCB7C435,
32'hBD9E30B8,
32'hBD9103E1,
32'hBE8B1FE5,
32'hBDFE53DD,
32'h3E723608,
32'hBC551372,
32'hBD8511A7,
32'h3E05F680,
32'hBF27F175,
32'h3E6D20CF,
32'h3DFE7D27,
32'hBE926B34,
32'hBE46C115,
32'h3D5A7103,
32'h3D8C1359,
32'h5DC5E11A,
32'hBD94B9DF,
32'h3E2AE28F,
32'hBE94BB38,
32'h3DDCE02D,
32'h3D762ECD,
32'h3D18B243,
32'hBF8148D9,
32'h3E6148CD,
32'h3CB11495,
32'hBE8BCB9D,
32'hBDA02DF1,
32'h3D7F550F,
32'h3E2D10DA,
32'hBDA9CBBB,
32'h3CA28B20,
32'hBEA6FE3B,
32'h3CA9CC16,
32'hBED6AD42,
32'h3E419D8E,
32'h1DC423D6,
32'h5DC03E46,
32'h3E9239A8,
32'hBD919A9C,
32'h3E62DB0F,
32'h3E4F4DFF,
32'h3DA17800,
32'h3D85A699,
32'h3E724364,
32'hBE16BB8A,
32'h3D5470AD,
32'hBE26891B,
32'h3F1A1C58,
32'h3E0870BE,
32'hBEBD1829,
32'h3D22CFC0,
32'h5DF6DF00,
32'hBED5819D,
32'h3D964AA2,
32'hBEABEE9C,
32'hBE85E2C0,
32'h3E077A5F,
32'hBC8DD3F7,
32'hBEB14BC2,
32'hBDE64600,
32'hBC5B391B,
32'hBDDB7CDA,
32'h3CD8CF25,
32'hBEA9D215,
32'h3EBF28E1,
32'hBE69F0B0,
32'h3EC41204,
32'h3F009284,
32'h3EC6329C,
32'h3DF600E3,
32'h3F02DA13,
32'hBD907E9B,
32'h3D2B39D2,
32'hBD8E5508,
32'h5DEA8AF1,
32'h3DAB59B6,
32'hBDBA4726,
32'h3DD3D3A4,
32'h3E9805E7,
32'hBEE9F22B,
32'h2EC49F24,
32'h3E2F2E77,
32'hBE25A061,
32'h3E962613,
32'h3E050D64,
32'hBE2B0484,
32'hBE0A428B,
32'h3DA94964,
32'hBF0A3A78,
32'hBD722F38,
32'h0ECE7DC7,
32'hBE220296,
32'h5DDD3247,
32'hBDF54E5B,
32'h3E11446B,
32'h3E4E867F,
32'h3E6B59FD,
32'h3E3B4278,
32'hBDAFFEBE,
32'h3DACDBCE,
32'h3DC83BD8,
32'hBE87DF4F,
32'h3E160077,
32'h3D98E9AF,
32'hBE67D802,
32'hBE874303,
32'hBEF36C3B,
32'hBE4B15FC,
32'h3D5237F0,
32'hBE8E7F67,
32'h3E859EF2,
32'h3D05B35C,
32'hBE906063,
32'h3EDF6AF9,
32'h3CC561D5,
32'h3C576C2A,
32'h1CC15CB,
32'hBC5A4145,
32'h3EFA0242,
32'hBC82ECCD,
32'h3DA692DD,
32'h3D80D709,
32'hBE4397FA,
32'hBDA5E2A7,
32'h3C988870,
32'hBF5373E2,
32'h3F0E5DC9,
32'h3F01628E,
32'h3E4358CD,
32'h3EA10221,
32'hBD8B84CB,
32'h3E4FBB75,
32'hBE8C3DAC,
32'hBD800C43,
32'h3E3D7BFA,
32'hBED2E933,
32'hBF70776D,
32'hBE838414,
32'h3E266159,
32'hBEA61181,
32'hBE4325A5,
32'hBE1ACC1C,
32'hBDA66A6C,
32'h3E2C34FE,
32'hBE1A73AD,
32'hBDDF16A9,
32'hBC28E44C,
32'h3D2BE23F,
32'h3D9E3F60,
32'h3C41DE82,
32'h1751F755,
32'h3EBE161E,
32'hBE9258B6,
32'hBDA8F5AF,
32'h3E1C4C54,
32'hBFFC4092,
32'h3E23A582,
32'h3E83C9ED,
32'hBD7CB84D,
32'h3ECC3556,
32'h3E919343,
32'h3EE398E5,
32'hBDCB519C,
32'hBD98DA24,
32'hBF3C2B52,
32'h3E327FEE,
32'hBFE1CC48,
32'hBDC2B0A4,
32'h3DED5CC4,
32'hBDBAB5F3,
32'h3E0899AD,
32'h3E06E832,
32'h3E2151BB,
32'hBD651382,
32'hBD1BD180,
32'hBDE98058,
32'hBE310FED,
32'hBE8A8887,
32'hBF0B929C,
32'h3D04E26A,
32'hBD1909A6,
32'h3E9970FE,
32'hBE9CB74E,
32'hBE8666FB,
32'hBC3E5684,
32'hBFB8487E,
32'h3E93078D,
32'h3E71AA53,
32'hBD609AE2,
32'hBC96BB0F,
32'h3E94DD38,
32'h3E9E9768,
32'hBDB0EB0C,
32'h3F142CC4,
32'hBDCB795A,
32'hBCED9A5B,
32'hC01A34C4,
32'h3DB879E5,
32'hBE12A5E8,
32'h3EB2C86A,
32'hBDE5803C,
32'h3DDBC934,
32'h3E91392F,
32'h3F0586F1,
32'h3E97640C,
32'h3D80A5C0,
32'h5DE8B82C,
32'hBD425F48,
32'hBEF6E2C0,
32'hBD21C098,
32'h3D0C77ED,
32'h3EBDA570,
32'h3DE8293A,
32'hBE888B8E,
32'h3D09FC2F,
32'hBF76F138,
32'h3E6C9202,
32'h3D4E4820,
32'hBE88C699,
32'h3E6DF2E2,
32'h3CF61F71,
32'h3F652767,
32'h3E89AA8A,
32'h3EB49B4B,
32'hBE1BED41,
32'hBEE8CA5B,
32'hBFDB47AB,
32'hBC46387C,
32'h3EAD000F,
32'hBE61821B,
32'h3F23119E,
32'hBE40A941,
32'h3E6408F5,
32'h3E1CC2A9,
32'hBECB542C,
32'h3E58AD15,
32'h3E89E504,
32'hBD48DD48,
32'hBEDAEDF0,
32'hBD8A3B64,
32'hBD5B839E,
32'h3ED970B1,
32'hBCA3E7CD,
32'hBDDF92F4,
32'hBD8BECE8,
32'hBF6000A1,
32'hBE3A854C,
32'hBC6E9C07,
32'hBE3919B6,
32'h3E2407F4,
32'h3E7F9541,
32'h3D0545F7,
32'h3EB904C9,
32'h3E6D8622,
32'h3ECEEE08,
32'hBE7BEDC9,
32'hC013C1BC,
32'h3D22DC87,
32'hBE139C3C,
32'h3F62E2D8,
32'h3F13846C,
32'hBE9AFBEA,
32'h3F05A06C,
32'hBEE66521,
32'hBE560DE0,
32'h3F4DA9C1,
32'hBF0A078B,
32'h3D83E7C6,
32'hBEDE9FB5,
32'h3D6E6A6B,
32'h1DF81A62,
32'h3F08F4F7,
32'h3E1A645E,
32'h3E253AA4,
32'h3EB13B15,
32'hBED76A3B,
32'hBE2303FC,
32'hBF292DD6,
32'hBECEF3F6,
32'hBF22F4DB,
32'h3D1CB161,
32'hBF844E05,
32'h3F0EC2CA,
32'h3F45D72B,
32'hBED668BA,
32'hBEE627F0,
32'hBF43EDAA,
32'h3E0D42D3,
32'hBEBA4796,
32'h3F6AB6FE,
32'h3F21100F,
32'h3D7ADB78,
32'h3EC01420,
32'h3F939004,
32'hBED59F4A,
32'h3F9C274A,
32'hBD29BC0C,
32'h3F02930E,
32'h3E33251C,
32'hBCF60BCE,
32'h3C993AA5,
32'h3EA20B66,
32'hBCCB3B4A,
32'hBE93F656,
32'h3EC06E3B,
32'hBE6B0556,
32'h3E2B2B06,
32'h3EB775A9,
32'h3F14EFA6,
32'h3E303FE2,
32'hBEFBA22B,
32'hBF40720E,
32'h3E1A20D1,
32'h3EDC87B0,
32'h3EE6F1F6,
32'hBF0CF382,
32'hBC95F370,
32'h07580EE2,
32'hBEC46F7F,
32'hBF2E1C35,
32'h3D633BE1,
32'h3F4F9598,
32'hBEF0E0ED,
32'h3EF2CD85,
32'hBE9867C7,
32'h3F804612,
32'h3EF787EA,
32'h3F9013E3,
32'h3FAF1852,
32'hBDADE70C,
32'h3D6572D6,
32'h3E8BA786,
32'h3F2D9E3D,
32'h3E2E32B3,
32'hBD3200C5,
32'h3F6C13BD,
32'h3E435D65,
32'hBF6EB2BA,
32'h3ED37EE8,
32'hBF7E1FBC,
32'hBF269035,
32'hBEEA9E37,
32'hBEAF1651,
32'h3F613F3C,
32'h3D01DEDA,
32'h3EFE747E,
32'hBDB07A14,
32'h3F391D25,
32'hBE2124D5,
32'h3C7AF6AB,
32'hBD86144C,
32'h3EF290F4,
32'hBCFBF3D1,
32'hBC836DEA,
32'hBDA4082A,
32'h3ED008A8,
32'h3EAC1B44,
32'h3F005C7B,
32'h3E70DF1D,
32'h3DC08DD5,
32'hBCF4C277,
32'h3CA961F3,
32'h3F063B3D,
32'h3DE6B2C4,
32'hBA406F5,
32'h3F0D8E06,
32'h3D245806,
32'h075B60B9,
32'hBE22C76D,
32'hBE23C657,
32'hBE7234B9,
32'hBD194477,
32'hBECE2150,
32'h3EE8057B,
32'h3CEDF2E9,
32'h3EC33C25,
32'hBD80ECA2,
32'h3F0E6189,
32'hBEB9F6C1,
32'hBC08FD84,
32'h3D0DD7C5,
32'hBD1EA2D4,
32'h3D1DEF81,
32'hBDC96A62,
32'h3F20E338,
32'h3E35D511,
32'h3E2DFD70,
32'h3CBD05B1,
32'h3D40B383,
32'h3D270167,
32'hBD44883E,
32'h3C9A3FEE,
32'h3D786F47,
32'hBD1BE212,
32'hBEA8D222,
32'h5DD16B84,
32'h3D8BECE3,
32'hBE5C2374,
32'hBDA06A57,
32'hBDBD54A8,
32'h3F1645D4,
32'h3DC0AB1F,
32'h3DBB3F47,
32'hBE06F9BE,
32'h5DCBDB57,
32'h3F67B20D,
32'h3DC81E10,
32'h3DC336CB,
32'hBC88BBCE,
32'h3D23DA98,
32'h5DFB249E,
32'hBD270E65,
32'h3C8E6050,
32'h3D124866,
32'h3D3E5881,
32'hBD1DDC28,
32'h5DEF4BDD,
32'hBD064625,
32'hBCF34B09,
32'h3DC74847,
32'hBD9F4F77,
32'h3D082CF7,
32'hBE8C3E84,
32'hBD3A0BFB,
32'hBE7AABD2,
32'h3DA539A9,
32'h3D05C231,
32'hBD49C0D1,
32'h3D473275,
32'h3C2EAF3B,
32'h3E98E5FD,
32'h3D5C1298,
32'hBCD7C9DC,
32'h3E657F39,
32'hBD2C91D4,
32'h3DBC1788,
32'hBDA26197,
32'hBCA8BF6A,
32'h3D83F712,
32'h3EA4B489,
32'h3DD8A659,
32'h3E52649E,
32'hBDD45938,
32'hBCA49F8E,
32'hBDE28B26,
32'hBEA3D5CD,
32'hBDB67F07,
32'h3E16D7E1,
32'hBDA9D843,
32'h1DC317B0,
32'h3D9C065B,
32'h3D1D573E,
32'hBE8A8629,
32'hBE732FBE,
32'hBF1595EF,
32'h3F1D854A,
32'h3EF21AF4,
32'hBF73AF18,
32'h3F96D376,
32'hBE217FC4,
32'hBE91A11B,
32'h3D580ADE,
32'hBE34D990,
32'hBCCACF7A,
32'h3F35F14E,
32'h3E201D7D,
32'h3CC9933C,
32'hBF19F7E9,
32'h3F9589CF,
32'h3E40E53C,
32'h3F166EFD,
32'hBEF592BA,
32'hBF6399D9,
32'h3F14E703,
32'hBDB17266,
32'h3E91F26E,
32'h1DE96C62,
32'hBEC609D3,
32'hBE3A95EF,
32'hBD049087,
32'h3CA3222B,
32'hBEE20075,
32'h3F351ADC,
32'hBE106D2E,
32'h3F7D5C18,
32'h3DF5F105,
32'hBE3C146E,
32'hBDA421CA,
32'hBDFD655E,
32'hBE55CA12,
32'hBF6674C6,
32'hBEE347D3,
32'h3DAE2EEA,
32'h3D2F2A43,
32'h3F8B9502,
32'h3E8CB7CA,
32'h3E7B2A89,
32'h3DA23B96,
32'h3ED73865,
32'h3EA4B24B,
32'h3E54DF39,
32'h3C96270A,
32'h3C0FBDF2,
32'h3F157C0B,
32'hBF0EC192,
32'h3DD14E26,
32'h3E06F6C5,
32'hBEDFEC07,
32'h3F1F70EA,
32'hBCF6DD5B,
32'h3DC683A3,
32'h3DF812CE,
32'h3F4EB64B,
32'hBE9D967D,
32'h3EF69095,
32'hBEE4DBEF,
32'h3F0E3684,
32'h3EE958FB,
32'hBD773A2C,
32'h3E7B48FB,
32'hBDB4C809,
32'hBE2D3BC5,
32'h3E3DBBFE,
32'hBF20D3E3,
32'h3ED88367,
32'hBEF97EB5,
32'h3E089F06,
32'h3F4CBA8E,
32'h3F0460E1,
32'hBE8B1D45,
32'hBE592BA2,
32'hBEC9134A,
32'h3ED97A0F,
32'hBE02B633,
32'hBF38EF44,
32'hBEE379AE,
32'h3EBA16F3,
32'hBF8B4270,
32'hBEB1A42A,
32'hBCBD670B,
32'h3DBD010B,
32'h3E183772,
32'h3D35CBC1,
32'hBF6DF8AE,
32'h3E136C17,
32'hBEF9B418,
32'h3CEA3944,
32'h1DFDD67B,
32'h3DF1AC42,
32'h3DEF0421,
32'h3E420894,
32'hBE30E540,
32'h3E2DBCCA,
32'h3D151EFD,
32'h3F2F438B,
32'hBC2A66A4,
32'h3EDE5105,
32'h3F5978BB,
32'h3F3B2C63,
32'hBEE7D7BF,
32'h3EBD408C,
32'hBF7408AB,
32'h3EA8A6AB,
32'hBC96D453,
32'hBEF52412,
32'h3D931B0B,
32'hBC14EB88,
32'hBF91925C,
32'hBF57D3AE,
32'hBD8826A7,
32'h3C81D728,
32'h3E4B5F25,
32'h3F3F845F,
32'hBE29A908,
32'hBE435668,
32'hBF6631E3,
32'h3E998C3D,
32'h3D7A6763,
32'h3E3927BE,
32'hBE3E8B52,
32'h3E6DF66A,
32'h3ECF9F7F,
32'h3E942FC1,
32'h5DE52688,
32'hBDDE4847,
32'h3DE574E4,
32'h3EA62122,
32'h3EDC8765,
32'h3E62352C,
32'hBCD84798,
32'h3E459AFD,
32'hBFB0426C,
32'h3F4B9567,
32'h3E89D1B6,
32'hBF3A853B,
32'hBEA84418,
32'hBE71AA04,
32'hBEFF5CC7,
32'hBEB679B9,
32'hBD95FC78,
32'hBDB159D5,
32'h3EAF684C,
32'h3E0898FA,
32'hBF0F427A,
32'h3E1204EF,
32'hBE07FB81,
32'h3C648DE6,
32'hBE07FCB4,
32'hBE0C00CC,
32'h3E3FDC3F,
32'h3D5263A7,
32'h3EEDC8CA,
32'h3E9926D8,
32'hBD841DA9,
32'hBC1B1558,
32'hBD7E09AE,
32'h1DD3EF44,
32'h3DB7133C,
32'h3F043C29,
32'h3E985934,
32'hBCB1E592,
32'hC028560F,
32'h3E8630C7,
32'hBDB9AEF2,
32'hBF133DD8,
32'hBF368B81,
32'hBF12AA75,
32'hBE9FEF79,
32'h3DCB8A11,
32'hBDB039BD,
32'h3D0D684F,
32'h3EC33FA6,
32'h3EF74B6A,
32'hBE3FC134,
32'hBDC79683,
32'h3E20DB39,
32'h3DC2AB30,
32'h3E5F362E,
32'h3E65F1FE,
32'h3E6387E4,
32'h3DDDD142,
32'h3ED46842,
32'h3E8A2AE4,
32'hBE1452F1,
32'hBF3204B2,
32'hBE344421,
32'h3E2452CF,
32'hBDA4F332,
32'h3EF1A52B,
32'h3E74CA2B,
32'h3E894BC0,
32'hBFBBFF70,
32'h3EBEC8B5,
32'h3D84AAD6,
32'hBE27141D,
32'hBEFF263F,
32'hBE9CC292,
32'hBCDF2DCC,
32'h3F1A1C6C,
32'hBE0A0827,
32'h3DA1B9FD,
32'h3E954649,
32'h3F483135,
32'h3E2320C4,
32'hBC05C73A,
32'h3F045B92,
32'h0ED1FC54,
32'h3CA3330E,
32'h3E06965B,
32'hBD268831,
32'hBD319A2B,
32'h3EEEC4CA,
32'h3D73C2E2,
32'h3E51F71C,
32'hBF6120F9,
32'hBCDCA35C,
32'h3D9CC383,
32'hBE0088E9,
32'h3EDD5102,
32'hBD6779CA,
32'h3F29A23B,
32'hBEE4E6BC,
32'h3E3A6531,
32'hBE509D66,
32'hBD9A1B8E,
32'hBE6CF43D,
32'hBE865167,
32'h3E0076F8,
32'hBF3C740B,
32'hBC4E4BE7,
32'hBD8A2041,
32'h3DFE9ED2,
32'h3E8CA529,
32'h3E261F8C,
32'h3D1D91CA,
32'h3ECC6AF4,
32'h3E7BD7EF,
32'h3E11331A,
32'h3E81C93B,
32'hBD6AC2E5,
32'hBD8F9FC3,
32'h3EA6801D,
32'h3DEEC8B1,
32'h3E1FB529,
32'hBF352FAB,
32'hBE7058F5,
32'h3E6F8F6E,
32'h3D4AFFAD,
32'h3F2B2DA1,
32'h3EACC3C8,
32'h3E199745,
32'h3E1E1ED9,
32'h3E56F91D,
32'hBDF6F5DF,
32'hBEB83C5E,
32'hBE14538E,
32'hBEE1C08F,
32'h3E098CDC,
32'h3E704D49,
32'hBC888500,
32'h3D236E55,
32'h3EB1E8AA,
32'h3DFCC951,
32'h3F160967,
32'h3CBE012F,
32'h3DEA88E5,
32'hBCCD08D5,
32'h3DC4D3C4,
32'h3DDA5E5C,
32'h3DECF4AD,
32'hBDD06B28,
32'h3D43D673,
32'hBE03C904,
32'h3E45425B,
32'hBF2A698A,
32'h3D535D27,
32'h1DE51F7E,
32'h3CAF70BB,
32'h3EB9BFD4,
32'h3E4EAD00,
32'hC0101D4B,
32'hBD40E736,
32'hBE051189,
32'hBDB21BAE,
32'h3CBD4E62,
32'h3D3DCAFC,
32'hBEB62766,
32'h3EB096EC,
32'h3E16D428,
32'hBDC273B6,
32'h1DDAF5D1,
32'h3CABDDFC,
32'h5CF9FA2,
32'h3ED1B5AC,
32'h07529ED9,
32'hBDAFF184,
32'hBE79992A,
32'hBEA9A592,
32'h3E97AC91,
32'hBDFF0216,
32'hBE87D296,
32'h3E78C5F1,
32'h3C95AFAB,
32'h3E94EE07,
32'hBF534E9A,
32'h3CA4577D,
32'hBE2CC80D,
32'hBE40530E,
32'h3CC44E67,
32'h3DE77DAA,
32'hBFF4E717,
32'hBE68DF31,
32'hBF03DC4E,
32'hBE215D2E,
32'h3DD7E4C4,
32'h3E75780F,
32'hBEAC4722,
32'h3E945892,
32'h3E32783B,
32'h2EDC1E2F,
32'hBCADD5AD,
32'hBEC9E219,
32'h3D9602DB,
32'h3E49BC81,
32'h3E61B158,
32'h3D9D22E7,
32'h07585661,
32'hBE9C84DD,
32'h3C38702B,
32'h3DA8B323,
32'hBD314F19,
32'hBDCD7FC8,
32'hBD9B2681,
32'h3E993EE2,
32'hBE3CD2A4,
32'h3E04E1E7,
32'hBD866CB9,
32'hBE7534F3,
32'hBE0EC51A,
32'hBE7B9ACD,
32'hBF0B594D,
32'hBDB7EBE1,
32'hBF834D94,
32'h3E8B0D98,
32'hBD0CD50E,
32'h3EAD7D32,
32'hBE65FE50,
32'h3CAB69A0,
32'h3D884D23,
32'h3D972663,
32'hBCA7C4B2,
32'hBDB9FB08,
32'h3E1BC15A,
32'h3C692B48,
32'h3EB1E3A2,
32'hBE0E3198,
32'hBD8FE3D7,
32'h3DB56E9C,
32'hBEADAFB9,
32'h3E26A08D,
32'h3E5FA462,
32'hBEFD8B0F,
32'h3D9EDCE4,
32'h3CA11025,
32'h3DCD7350,
32'h3E5E601B,
32'hBDD32D53,
32'hBE80BBE9,
32'h3D3CD226,
32'hBE552338,
32'h3DC45A82,
32'hBC9023A3,
32'hBF7F6DC6,
32'h3E6F202B,
32'hBD98E162,
32'h3D5265AE,
32'hBEA772BA,
32'hBC9F628B,
32'hBEBC9A40,
32'hBC9B031E,
32'h3D6D8729,
32'hBE031283,
32'hBE7C195D,
32'hBE34AD22,
32'h3E91E4DB,
32'hBE57CAB0,
32'hBDEDC4C2,
32'h3E9434B4,
32'hBEE8F1F3,
32'h3F05F2AB,
32'h3EA4F1B8,
32'hBE4F4094,
32'h1DE52C44,
32'h3DC83AC0,
32'h5DDB1B40,
32'h3E0AFEAB,
32'hBE183CBB,
32'h3D8D8871,
32'h3DB6E304,
32'h3DA94372,
32'hBE263413,
32'h3DCA2B91,
32'hBEBAD7A5,
32'hBE79A6E5,
32'hBDDAE40D,
32'hBE963FB8,
32'hBE59D322,
32'h3EBCE422,
32'h3EB502FC,
32'hBDBEB9F7,
32'hBD333660,
32'hBD646A07,
32'h3D4E84AC,
32'hBA02234,
32'h3E051553,
32'h3EB05A7A,
32'h3CE68403,
32'h3EBB00D1,
32'h3CA020EA,
32'h3E783A7B,
32'hBD1096D2,
32'h3E44921B,
32'hBD08E42D,
32'h3C584EA6,
32'hBDA8F9A6,
32'hBCBB23AD,
32'hBDA8C21B,
32'h3EE1A86B,
32'h3E8256EE,
32'hBD9AA48D,
32'h3DDD6B67,
32'h3DFDA0E7,
32'hBF0F1F59,
32'h3E671573,
32'hBE8C8751,
32'hBD54AC7C,
32'h3DD568C1,
32'h3E032F5A,
32'hBF1D9ED8,
32'h3D54C6C2,
32'h3D5DF7D2,
32'hBE155D84,
32'h3E2DC3C6,
32'h3DD2FE5E,
32'h3DB6E17B,
32'hBF0807F8,
32'h3DB3DE2B,
32'h3ECCFE6A,
32'h3E352B69,
32'h3E5D03BC,
32'h3E0709EA,
32'h3E1CC432,
32'hBC97C0D2,
32'h3DF5A12B,
32'h3EF16C64,
32'hBD7EF6E7,
32'h3D1D1F52,
32'hBC7CF8A6,
32'h3EC3BA1A,
32'hBEF08A4D,
32'h3E0F956C,
32'h3DAB824C,
32'hBD8C0E18,
32'h3E217291,
32'h3E7397F1,
32'hBE0BF29D,
32'h3E0F0F47,
32'hBDDA1751,
32'hBF55731F,
32'hBD323E1E,
32'hBD60F372,
32'hBE75DD8A,
32'hBE80BA1E,
32'hBE1D4E23,
32'hBD058D0C,
32'hBFEC0D46,
32'h3DAFA7E6,
32'h3E89DB22,
32'hBC92B590,
32'h3E77620A,
32'h3E225F20,
32'hBD6353D4,
32'h3DC68CB4,
32'h3E55AB89,
32'h3EADC9FB,
32'hBECF8405,
32'hBCBA3B28,
32'hBE81ACF1,
32'hBE674468,
32'hBF1F68E4,
32'h3E8831A5,
32'h3D83CE73,
32'hBE9D7FDF,
32'hBCBD28E9,
32'hBC6D0FA2,
32'h3D9C527D,
32'h3DB6E798,
32'h3E75AC8A,
32'hBE49DE6A,
32'hBD95AA6F,
32'h07583626,
32'h3E9E3F62,
32'h3E47498C,
32'h3E042BD9,
32'h1DFECCD7,
32'hC0199774,
32'hBCA36982,
32'h3E98BC97,
32'h2EC9438C,
32'h3E904F18,
32'h3D0F163A,
32'h3E8CD883,
32'h3E09F34E,
32'h3E8D500E,
32'h3F152299,
32'hBDACE171,
32'hBEEC5884,
32'h3C60EE05,
32'hBE1EFA93,
32'hBF401F96,
32'hBD652DD2,
32'hBE8A7277,
32'hBDF0D983,
32'h3D865F47,
32'h3C017F19,
32'h3EC8C1DF,
32'h3CA09679,
32'h3F173B87,
32'hBF1A7BF6,
32'h3C96507E,
32'hBC115E54,
32'h3E8A746B,
32'hBE1EBD85,
32'h3E25FF16,
32'h5DD8F0B3,
32'hC0121593,
32'hBE097FC2,
32'h3F1132FA,
32'h3E8B33C8,
32'h3DFE9742,
32'h3E509A9C,
32'h3EA2816F,
32'h3E4C0EDF,
32'hBCB70B94,
32'h3DFF3548,
32'h3E064B56,
32'hBF71447A,
32'hBD9DCB0B,
32'h3E85861A,
32'h3E88DC25,
32'h3D86B725,
32'hBC47EE8E,
32'h3E2EA0D2,
32'h3DAD56E0,
32'hBE0013B5,
32'h3DC966E6,
32'hBE067DF0,
32'h3E13ED4B,
32'hBE4DAAA7,
32'hBD16A98A,
32'hBD7DCC50,
32'h3D56C16E,
32'h3E774F5E,
32'hBD404E8A,
32'hBEA42348,
32'hBF7F3204,
32'h3CB981B6,
32'h3EF7E5B4,
32'hBD7236AC,
32'h3E9A41E2,
32'h3DE99C53,
32'h3DA1D400,
32'h0ECE6D54,
32'h3F0EC16A,
32'h3F44FDE7,
32'h3C891E4A,
32'hBF8421E2,
32'hBE4DB33B,
32'h3E2EE0A3,
32'h3EF5057B,
32'h3D914BB7,
32'hBE404C65,
32'h3D23AE23,
32'h3E7E6CCB,
32'h3E7C44E8,
32'h3D9F06B6,
32'h3DC66FA8,
32'h3DBBD9E8,
32'hBDEFB566,
32'hBD91C81F,
32'hBD9E36BB,
32'h3E59C873,
32'hBD5D75CA,
32'hBCDBAB4C,
32'hBD07D316,
32'hBF19DAD7,
32'h3DD394E9,
32'h3EA2589C,
32'h3DB19722,
32'h3EAF3376,
32'h3E068E3C,
32'h3F478A8D,
32'h3E8215B1,
32'h3F40D357,
32'h3DDF5E99,
32'hBEB22B79,
32'hC00729BB,
32'hBE968BF4,
32'h3EA958CD,
32'h3E56CF72,
32'hBDC9CD23,
32'hBE9CD08B,
32'h3E43A60A,
32'h3E89DE27,
32'h3EEE7798,
32'h3EDF99FF,
32'h3E468CAA,
32'h3ED98A5E,
32'hBDD548E5,
32'hBDE56412,
32'h3DCEAA5B,
32'h3DB28F62,
32'hBEA877EE,
32'hBE14CC94,
32'h3D9FCB3C,
32'hBDE1A9C6,
32'hBE7E2411,
32'hBCCA2394,
32'h3CE6658C,
32'h3E30BBB1,
32'hBD0DCD69,
32'hBE7D9104,
32'h3F06C5C1,
32'h3EEE9D74,
32'h3EBF4582,
32'hBEAFB315,
32'hBFD58B74,
32'hBE03578D,
32'h3E9D3206,
32'h3F41E99B,
32'hBF1A318F,
32'h175B484A,
32'h3F314EE7,
32'h3E41D4A7,
32'hBE285DFC,
32'h3F4791E6,
32'h3EB457E8,
32'h3EE9A24D,
32'hBC659964,
32'hBDDE5D85,
32'h3C08756F,
32'h3E854FC0,
32'h5DE69F0F,
32'h3EEE07FF,
32'hBD957251,
32'h3F111469,
32'hBE593AF3,
32'hBEE2C129,
32'hBF07816C,
32'hBF099366,
32'h3E169150,
32'hBF645634,
32'h3F105C2B,
32'h3F625AA1,
32'hBD36BFAA,
32'h3EDF25A0,
32'hBFC2B78E,
32'h3EA0BCFE,
32'hBECDF53C,
32'h3EB5052E,
32'h3EC0CFA9,
32'h3E3C1C53,
32'hBD7DEB03,
32'h3E9FE736,
32'hBF298088,
32'h3FA52BC8,
32'h3E5DC395,
32'h3F210E88,
32'h3ED8E74C,
32'hBDA5EDB8,
32'h3DC7334A,
32'h3EEF8164,
32'h3E7531B2,
32'h3E8BF5D9,
32'h3E2B3118,
32'h3F075C60,
32'hBD05ABC6,
32'hBF3B4AED,
32'h3E8C521C,
32'hBE90AF39,
32'hBE348494,
32'hBF5AE13B,
32'h3F712E90,
32'h3E128A19,
32'h3DA5F14F,
32'h3E2B6573,
32'hBEBA510D,
32'h3F012DE4,
32'h3DDC01FE,
32'hBF484306,
32'hBD124E7C,
32'h3F3B1C78,
32'hBF8682C8,
32'h3D6F69F5,
32'hBEDA90DC,
32'h3F7C690A,
32'h3EFE4650,
32'h3F6D17B5,
32'h3F80D62C,
32'h3D020AEA,
32'h3D99F864,
32'h3E289B91,
32'h3F3E397D,
32'h3E5B15FD,
32'hBE8226A3,
32'h3FB4CF42,
32'hBF2190ED,
32'hBFA1EE2F,
32'h3D259F16,
32'hBEEA2667,
32'hBF545009,
32'hBF7A8503,
32'h3EBF0D6C,
32'h3F371719,
32'h3ED6554D,
32'hBE9B85DC,
32'hBDD873E2,
32'h3FA04AB2,
32'h3E767BE5,
32'hBD62E09D,
32'h3C8E22A2,
32'h3F691764,
32'hBECD2646,
32'hBE0CDEB2,
32'hBDC43249,
32'h3FA21DDF,
32'h3F2E390F,
32'h3FAB2CCD,
32'h3DE8F86D,
32'h3D368DAF,
32'h175E2CB5,
32'hBEA290AC,
32'h3F38105E,
32'h3DA52236,
32'hBD9109EE,
32'h3F49BBCA,
32'h3D11E4F6,
32'hBC75FFD8,
32'hBECC67BC,
32'hBD844CBE,
32'hBF042F93,
32'hBE594118,
32'hBFA11B7C,
32'h3EF0F57C,
32'h175FAC76,
32'h3F98809A,
32'hBD76EE07,
32'h3F30D929,
32'hBF4DCCB1,
32'hBD130081,
32'h3D0538A1,
32'hBD98ACBF,
32'h3C807815,
32'h3D0419A9,
32'hBD0492FA,
32'hBD9882EA,
32'h3DA0EF2A,
32'hBD16B172,
32'h3C61E506,
32'h5DD120DE,
32'hBD185BF7,
32'h3CF14A65,
32'h3C9409E1,
32'h3DB2EA7D,
32'h3C9E0AC2,
32'h3CD7056C,
32'h3D53B6D9,
32'hBDB3547D,
32'hBCAC49B1,
32'hBC94AB99,
32'h3E2F398D,
32'hBC356AC3,
32'h07586035,
32'h1DE65B64,
32'h3CEC44AA,
32'h3DB73EA3,
32'hBCCE86B8,
32'h3DDCB5B5,
32'h3DD27C12,
32'h3D737604,
32'hBC2D7550,
32'hBD6FF13C,
32'hBD84DEA4,
32'h3D84BCEF,
32'hBCA833ED,
32'h3F0544A5,
32'h3F39C3D9,
32'h3DC2F174,
32'hBD8FCB01,
32'h3D69EDED,
32'hBD5AC0EB,
32'hBD6FBC3D,
32'hBEC26C60,
32'hBDD0459B,
32'hBE2C70B4,
32'hBD4DF163,
32'hBD049AD2,
32'hBD34118D,
32'hBDE4A120,
32'h5DFDD017,
32'h3E9C1D50,
32'hBCD7A11D,
32'hBF6AD66F,
32'h3F767006,
32'hBD9ACAF4,
32'h3F0B7F2B,
32'hBC726C30,
32'h3E98F60F,
32'h3D042115,
32'h3EC9E751,
32'h3E10CC84,
32'h3FB7F199,
32'hBEB41309,
32'hBDC6A935,
32'h3F115502,
32'h3F14B748,
32'h3EEC5EEA,
32'hBCE8EBA3,
32'hBE283504,
32'hBD4DFEF0,
32'h3CA5E64C,
32'hBDEA357C,
32'hBEA18281,
32'h3EC65FFA,
32'hBE8DCA27,
32'h3F1C7380,
32'hBDF7556A,
32'hBF8FB958,
32'h3F2FB16F,
32'hBE8F2EFD,
32'hBEB6F132,
32'hBD8BF8EE,
32'hBF8130F2,
32'h3F4E7EFE,
32'h3EFB32E6,
32'h3F554F68,
32'h3E9F8600,
32'hBEF337AF,
32'h3F64D509,
32'hBD82866C,
32'h3ECBEE7B,
32'hBE2D305C,
32'hBFDAA800,
32'h3F0008B0,
32'h3D31CC50,
32'hBEB8BD1D,
32'hBE2F2AEE,
32'h3ED5B31F,
32'h3E4E8A3A,
32'hBDB425BF,
32'h3D5AE331,
32'h3CE1DE68,
32'hBD91CF40,
32'hBED6072E,
32'h3F535DB8,
32'hBE7499F4,
32'hBEA16D4E,
32'hBF0E7DA8,
32'h3DA09943,
32'hBEEAD298,
32'h3D9B22BE,
32'hBEBE59FC,
32'hBE3F7459,
32'h3F5A47B9,
32'h3F1E27CC,
32'h3F342777,
32'h3E5B9F0D,
32'hBCEDE8CF,
32'h3E80556E,
32'hBF427342,
32'h3F6AEE88,
32'hBF95B7C7,
32'h3F0459E5,
32'h3C648127,
32'hBDA8A83A,
32'hBDAFE9AA,
32'h3ED21B68,
32'h3E28A09A,
32'hBD8C4CD2,
32'hBDADCCFF,
32'h1DC53A5A,
32'h3E2D3895,
32'h3EBD9494,
32'hBF2D00B9,
32'hBD70C021,
32'h3E012A0A,
32'hBEBAF387,
32'h3CADE154,
32'hBEA7C7FB,
32'h3E919152,
32'hBE0D66FB,
32'hBF0709B4,
32'h3D1B0F51,
32'h3F62CB02,
32'hBDF262E8,
32'hBEC12F46,
32'hBCB5E68A,
32'h3F13CDDA,
32'hBE9B5914,
32'hBF15669B,
32'h3CD30806,
32'hBF8D856B,
32'h3E9FB7C5,
32'h3E895B59,
32'h3DE7DD9B,
32'hBEAE9C10,
32'hBD6D6A59,
32'hBE0A30DE,
32'hBEB621AA,
32'hBD6FA094,
32'h3DDEB080,
32'h3DC0F4A8,
32'h3E60865F,
32'hBF26185E,
32'h3EA36414,
32'h3E7DCB7D,
32'hBE81C012,
32'hBDB7E6A0,
32'hBD90DD0D,
32'h3E266292,
32'h3DAEC923,
32'hBF5959E7,
32'h3E54D336,
32'h3D37F76A,
32'hBD9B68DD,
32'h3DC8BB1A,
32'h3F07FD76,
32'h3EFB54B7,
32'h3E859DA3,
32'hBEC3052A,
32'h3ED0F64E,
32'hBFCAB83D,
32'h3EEF0D4B,
32'h3D57C4DB,
32'hBF07D697,
32'hBEF243A2,
32'hBD161AAF,
32'h3EA9B28F,
32'h3F3DEB16,
32'hBCDD461A,
32'h3D08E381,
32'h3EDFAE72,
32'h3F0B53A3,
32'h3E99BADD,
32'h3E81C8CE,
32'h3F2B2937,
32'h3DBCBDF7,
32'h3DB08294,
32'h3E4715DF,
32'hBE3AFCDA,
32'hBDFE7CB2,
32'h3D9E0F99,
32'h3E9120D4,
32'h3E2F35C0,
32'h2EC806B4,
32'hBD8CA8C8,
32'h3E83D293,
32'h3DF7471A,
32'h3EB91955,
32'hBD2421F4,
32'h3EFF9A3F,
32'hC00ACA7D,
32'h3F30FE98,
32'h3E1BC526,
32'hBF54A1E4,
32'hBEF2E7D1,
32'hBEE93379,
32'h3E03DEA7,
32'h3D903365,
32'hBD45CF72,
32'hBC4EB299,
32'h3DBFD53F,
32'h3DFA0C25,
32'h3E1A1200,
32'h3E7E10D0,
32'h3F1F9468,
32'h3E600AD2,
32'h3EC5F750,
32'h3E858842,
32'h5DCBFE28,
32'hBD6C06AF,
32'h2EC46C40,
32'h3ECB3680,
32'h3E0BD31E,
32'h3E2829B5,
32'hBE0EC0C5,
32'hBDCBCFE6,
32'h2E59E91,
32'h3F1181AC,
32'h3E856E9B,
32'h3EA38F26,
32'hBFB204DF,
32'h3F121100,
32'h3D9BDCA9,
32'hBF9C7052,
32'hBF346334,
32'hBEF3A3DE,
32'hBE8BC503,
32'hBF2093EC,
32'h3CC04DA0,
32'h3D25E755,
32'h3E6ECF68,
32'hBDD318B4,
32'h3EAFE313,
32'h3E237971,
32'h3E4DCED2,
32'hBC84A6CA,
32'h3E8672A4,
32'h3ECFF562,
32'h3E48597A,
32'h3E0CF951,
32'h3E46FEFF,
32'h3EB444AB,
32'h3C934CB3,
32'hBE8B8622,
32'hBDE08511,
32'h3D062699,
32'hBEA9644A,
32'h3EE2F573,
32'hBDA759BA,
32'h3E8AADFE,
32'hBDAC3834,
32'h3F0853D3,
32'hBE2595D4,
32'hBF3D4975,
32'hBED7B610,
32'hBEE8569E,
32'h3D6F8F14,
32'hBD000E5F,
32'hBCF720E5,
32'h3D736F37,
32'h3E451840,
32'h3ECAF131,
32'h3EAD9307,
32'h3DA7000D,
32'h3E0859AD,
32'h3E66ADBA,
32'hBD8D4FBA,
32'h3EB0782A,
32'h3DB8AF89,
32'hBE390679,
32'h3E8CA6B7,
32'hBD74314A,
32'h3E656405,
32'hBF445EAC,
32'h3DE3AF1D,
32'h5DE9942C,
32'hBD7B61C1,
32'h3E955DD8,
32'hBEBD0531,
32'h3F4E5930,
32'h3EBDE234,
32'h3F0F86D3,
32'hBE0D5962,
32'hBEE1967D,
32'hBE5552C9,
32'hBF42CD07,
32'h3CD0905B,
32'hBE0DC103,
32'hBD8294F9,
32'hBCFE014A,
32'h3EECD336,
32'h3DC3B255,
32'h3EC57382,
32'h5DD01906,
32'h3DB3D2A1,
32'h3CCF4A77,
32'h3E4BA965,
32'h175081BA,
32'h1DED59C2,
32'h3D91B7FC,
32'h3E887595,
32'h3E4F29AD,
32'h3D8411CC,
32'hBF0AE5F9,
32'h3E137607,
32'h3E559CA0,
32'hBE571BAC,
32'h3E845A72,
32'h3E82F8B2,
32'hBF56B79F,
32'h5DF02EF6,
32'h3EDE7D8F,
32'hBEB1DEEB,
32'hBEA56D64,
32'hBF769F61,
32'hBF8C6B4C,
32'hBD9C6A83,
32'h3DAEBFF6,
32'hBD631C4A,
32'hBD9D2A3A,
32'h3EAA9259,
32'h3D94B51C,
32'h3EB1B3C9,
32'h3E245B2D,
32'h3E07E961,
32'hBE407BB0,
32'h3D0B78B6,
32'hBE9393AB,
32'hBDE76346,
32'h3E244F36,
32'h3DB78909,
32'h3E072C32,
32'h3C529F9D,
32'hBEC18CF5,
32'h3EE5119D,
32'h3E513CDD,
32'hBECFCAAC,
32'h3EAE41DB,
32'h3D66120C,
32'hC01130D3,
32'hBC64F265,
32'hBFA24246,
32'hBDEF0403,
32'hBE073AC3,
32'hBE55BE21,
32'hBF8F482D,
32'hBDECAE63,
32'hBE1D5028,
32'h2EC5C7E4,
32'hBD1A8DDF,
32'hBD3EDD9F,
32'hBD84F699,
32'h3DC9FD76,
32'h3E51BBDA,
32'h3E42371B,
32'h3D6F8581,
32'hBE127883,
32'hBE7F19C8,
32'h175D5E34,
32'h3CF6D5D0,
32'h3E322DC4,
32'h3E21AEB7,
32'h3F0B26B5,
32'h3DF8DB63,
32'h3E8401A3,
32'h3CD72E7A,
32'hBEC67143,
32'h3EADDBBD,
32'h3D2B5617,
32'hBF9CE3FE,
32'hBE089077,
32'hBF832C72,
32'h3E978BB2,
32'hBE12DAE2,
32'h3E6B5671,
32'hBF0A599D,
32'h5DC6DF81,
32'h3DAFAD0A,
32'hBD43FE30,
32'h1DF6CE9E,
32'hBE99D488,
32'h3D056C45,
32'h3E6AC1D9,
32'h3E649749,
32'hBDFC5D4D,
32'h1DD56CC6,
32'hBDF5D7E8,
32'hBD2CE6A5,
32'h3EE1CE0A,
32'h3E5B3CA5,
32'h3E6D20DD,
32'hBE6A9F70,
32'h3E6BE144,
32'hBE0CB663,
32'h3E83528A,
32'hBE44550C,
32'h3D87C002,
32'h3E334755,
32'hBE067737,
32'h3E20C595,
32'h3DA06E20,
32'hBFC31256,
32'h3E29FF9D,
32'h3E283F17,
32'hBE7A888A,
32'hBF197FC5,
32'h3EBEDED0,
32'h3DA6CC14,
32'hBDB135C7,
32'h17587761,
32'h3DE2CCC2,
32'h3D7E9773,
32'h3E42EA44,
32'h3E5978F3,
32'hBE80C113,
32'hBD55A5E2,
32'hBD2EF026,
32'hBE97228F,
32'h3E96BA68,
32'hBD0CD7B8,
32'hBEBEDD57,
32'hBDC3CF78,
32'h3D85BC4B,
32'hBDA2844E,
32'h3E10B10B,
32'hBE5C4D09,
32'h3E22277E,
32'h3CF9DF07,
32'h3DA3233A,
32'hBDB809F8,
32'hBE37A900,
32'hBEF0A6D5,
32'hBE2C4468,
32'hBE77A950,
32'hBE737962,
32'hBDB6A310,
32'h3EACD9E0,
32'hBC33DDBD,
32'h5DF1D5C6,
32'hBDAB9DDB,
32'hBD785356,
32'hBE407D15,
32'h3C94A953,
32'h3E6C5650,
32'hBE10F427,
32'h3E1F357D,
32'h3EBE5775,
32'hBE8968BD,
32'h3EB1D16C,
32'h3CCF03A2,
32'h3E1E705C,
32'hBDB583C7,
32'h3D7D9681,
32'hBDAB34FD,
32'h2ED8DA70,
32'h3DEB2B39,
32'h3ECBDE48,
32'h3EAD5219,
32'h3E599648,
32'hBEA89CB9,
32'h3DB077A5,
32'hBE513641,
32'hBDAAEE7C,
32'hBE074B95,
32'hBDB71A8A,
32'hBE813785,
32'h3E93D702,
32'h3E696BD1,
32'hBD118FBA,
32'hBD05B64C,
32'h3E354213,
32'h3E09B37F,
32'hBCCC133D,
32'h3E43DDA4,
32'h3E2C6831,
32'h3D1DA5DA,
32'h3E189CC1,
32'h3C328693,
32'h3EA523FD,
32'h3D84D03D,
32'h3DD295FB,
32'hBDBC3CAC,
32'hBDCA2EEE,
32'h3E1B09B1,
32'hBE1A0E58,
32'hBD18AACC,
32'h3E109C17,
32'h3EBAF9DF,
32'hBEC167A2,
32'h3E85F1E4,
32'h3E69F645,
32'hBE337732,
32'h3E1A6D60,
32'h3CA5BD08,
32'hBD43DF7E,
32'h3DD4ED90,
32'h3EC37A41,
32'hBF283DCB,
32'h5DEA7524,
32'h3C0670BC,
32'h3D78598C,
32'h3DE7E19E,
32'h2ECB448A,
32'hBCB5C2D3,
32'hBFCAA42C,
32'h3D190FC6,
32'h3E8B0F09,
32'h3D9855D3,
32'h3ED69D8E,
32'h3E721CB0,
32'h3DC35345,
32'h3D81F2EC,
32'hBC0103FA,
32'h3F02700D,
32'hBEA7D8D5,
32'hBE60820F,
32'h3E8AA194,
32'h3E2C053E,
32'hBD153D42,
32'hBD73799E,
32'hBD4BEFFA,
32'hBD72CC76,
32'hBD437ACE,
32'hBC51A9DC,
32'h3E1AF8D8,
32'h3DE7A234,
32'h3E6035F3,
32'hBF3DA2A7,
32'h0EC9B0E6,
32'hBDB92E5D,
32'h5DDB294D,
32'hBE8965EF,
32'h3E6E7F6D,
32'h3C81EB92,
32'hC0318ED2,
32'hBE27B2B9,
32'h3DCCA5B0,
32'h3C3BC396,
32'h3F060E5D,
32'h3EC5AB31,
32'h3CFBBAFB,
32'h3DC1AF37,
32'hBC33FD5C,
32'h3DE4595E,
32'hBE833DAC,
32'hBE2B3931,
32'h3DC53A49,
32'h3C7CF17E,
32'h3E1CF889,
32'hBD9AE662,
32'h3E9801D3,
32'hBE01B063,
32'hBC9FFE31,
32'hBE75D41E,
32'h3E7A832C,
32'h3E9B65CD,
32'h3EABDE42,
32'hBD4BE42A,
32'hBD31EFE1,
32'h3D7E59EE,
32'h3E321639,
32'h3E56EBEA,
32'hBCB9A41C,
32'hBDCA5082,
32'hC0168826,
32'h3C32036D,
32'h3E2A4F4E,
32'h3D869BB1,
32'h3E2A176B,
32'h3EC60AB2,
32'hBDA8AEAB,
32'hBD769DB9,
32'h3E892A04,
32'h3E2E17C5,
32'hBD0211C2,
32'h5DCF6105,
32'h3EB92AD4,
32'h3E6F7C3D,
32'hBC9D59B4,
32'hBE9CACEE,
32'hBE54D345,
32'h3E42EF9E,
32'h3E2AD4D8,
32'h3E77B479,
32'h3EBB87B8,
32'h3DA2F5DB,
32'h3E9DCD4B,
32'hBE0DD53A,
32'hBD513689,
32'hBD8BBD15,
32'h3EB80015,
32'h3CA368F8,
32'hBD87188E,
32'hBE251233,
32'hBF8EEC01,
32'hBED2A872,
32'h3E5A2EAF,
32'h3E2B99DF,
32'h3E65A6EC,
32'h3DF2A58D,
32'h3F019998,
32'h3E9E46F4,
32'h1DF39823,
32'hBE345E6C,
32'hBDD8825C,
32'hBE7D3A46,
32'h3E6D4F03,
32'h3F30B243,
32'h3EDADC2A,
32'hBD0F8D3A,
32'h3E7FBF34,
32'hBD8E21C9,
32'hBCB076E3,
32'h3D9D120D,
32'h3EE9C6A1,
32'h3DFDAD38,
32'h3E7E081B,
32'hBE2A224C,
32'hBCC07294,
32'hBCE5C338,
32'h3DF2E122,
32'h3E8E038C,
32'h3E3FD6F8,
32'hBDD39C25,
32'hBE821A49,
32'h07577268,
32'hBE2F7A08,
32'h3E964E23,
32'h3E9838F5,
32'h3E431DE5,
32'h3E487095,
32'hBCE6EE27,
32'h3E81BF56,
32'h3F302AFF,
32'h1DF37749,
32'hBF823A6E,
32'h3E5635A8,
32'h3F2B6BE5,
32'h3EBC1B70,
32'hBE88E337,
32'hBD3E8A84,
32'h1DE8BAA6,
32'h3EBC8431,
32'h3E9E2C05,
32'h3E6DC1BF,
32'h3F429921,
32'h3E545AE8,
32'hBD4BFF6F,
32'hBD5E8CE1,
32'h3CD21F8A,
32'h3E177C74,
32'h3E74EF01,
32'hBD50AD7F,
32'hBDAB1034,
32'hBE715BB8,
32'hBE23F6DB,
32'h3D9CB79B,
32'hBCF98C58,
32'hBE2A1419,
32'h3DEA77D5,
32'h3DCFEBCC,
32'hBD9D786F,
32'hBDE59197,
32'h3D9A3293,
32'h3DE39009,
32'hBFE4CD19,
32'h3E393976,
32'h3E6E10F0,
32'h1750931C,
32'hBF23DE2A,
32'h3EA675EB,
32'h0EC0A40D,
32'hBEC5F50C,
32'hBE9FB965,
32'h3F0FC152,
32'h3EC669DC,
32'h3EF02008,
32'h3EA10F36,
32'h3D723F22,
32'h3DE567BC,
32'h3D08BBA1,
32'h3E4BDE59,
32'hBE7DFC74,
32'hBDFF3674,
32'h3EA49E94,
32'hBEF37507,
32'h3DBCA8B9,
32'hBE38A077,
32'h3ECBE439,
32'h3D1B7B07,
32'hBF0E6A57,
32'h3DF2AFF9,
32'hBDE69527,
32'hBE0A374D,
32'h3DF20F74,
32'hBF7E5C9B,
32'h3DBCFC89,
32'hBDB473D7,
32'h3E5239C1,
32'hBF385AE3,
32'h3EEBA155,
32'h3D311B30,
32'hBEBA506C,
32'h3EA4342A,
32'h3F427444,
32'h075A04E2,
32'h3E388C21,
32'h3F8996CC,
32'h3D835F4D,
32'h3D9A1639,
32'hBDEC7536,
32'hBE90C587,
32'h3E700ECA,
32'hBDB59F68,
32'hBEAF0235,
32'h3E8BD2DA,
32'hBEE30E5A,
32'hBDE300DB,
32'h3EDA17AF,
32'h3E02157F,
32'h3E65D76F,
32'h3E2D0EFB,
32'h3E1D7DE2,
32'hBF839817,
32'h3F182816,
32'hBE9F42E8,
32'h3DAE72E8,
32'h3E487A0F,
32'hBE91482C,
32'hBF20085C,
32'h3FA0BCC7,
32'h3E59A8D5,
32'hBEF9C524,
32'hBF97F71F,
32'h3F97CA6A,
32'h3DA776D0,
32'h3F81C3E0,
32'h3F8ABEDE,
32'h2ECB00C5,
32'hBD73D2A4,
32'h3EE9BBA9,
32'h3EC0F8E3,
32'h3F4054F2,
32'hBEC4C7A0,
32'h3F38A597,
32'h3EB69BED,
32'hBFED9273,
32'h3E0819E7,
32'hBF17D74A,
32'hBEC4B893,
32'hBF656DCF,
32'h3F4043FC,
32'h3F93ED1D,
32'hBF0BD939,
32'hBD2198D3,
32'hBEAFF25C,
32'h3F1CBB0B,
32'h3E3C1B19,
32'h3EBDC7B7,
32'hBE04B08A,
32'h3F8F5B0F,
32'hBFA77FB7,
32'h3F697FA2,
32'hBE758ABD,
32'h3F42F42C,
32'h3E07DB17,
32'h3F58BDAE,
32'h3F258511,
32'h5DE6E9D8,
32'h3DF8256C,
32'hBD985666,
32'h3E8E5AA1,
32'h3E949C4D,
32'hBE07B41C,
32'h3FC9B688,
32'hBE3CFF8B,
32'hBF568922,
32'h3EA5E205,
32'hBEC18964,
32'hBEB3FFC3,
32'hBF6DE771,
32'h3EA4836D,
32'h3E98AA17,
32'h3F339026,
32'h3D8D4D88,
32'hBE92A795,
32'h3F42FDB5,
32'hBE9D43F2,
32'hBD07E245,
32'h3DC81F27,
32'h3F592AC7,
32'hBF11277F,
32'hBE37328D,
32'hBDC9FFFC,
32'h3FC4618A,
32'h3F2D9D23,
32'h3FA92441,
32'h3E19297B,
32'hBCE39205,
32'hBD849AF6,
32'hBE001965,
32'h3FA089CF,
32'h3D66DEE5,
32'hBEDF612E,
32'h3F4B292E,
32'h3D04F816,
32'hBED81220,
32'hBF082C35,
32'hBDEC2736,
32'hBECFB0D8,
32'hBD74BECD,
32'hBF7065C0,
32'h3F8239C0,
32'hBD2734C7,
32'h3FA1B464,
32'hBE19EADB,
32'h3F2863F7,
32'hBF94E2EA,
32'h3D64EF54,
32'hBC861A87,
32'h3D9601EE,
32'h3DAC722F,
32'hBD3C51D8,
32'h3D65A2CB,
32'h3D5528F4,
32'h3DCD6D30,
32'h5DF7E47D,
32'hBDE4CE74,
32'hBC3BE3E9,
32'hBDC20428,
32'hBD8BBAC5,
32'h3C286E59,
32'h3CA68CB1,
32'h3C7E0156,
32'h5DD15B0F,
32'h3CA5DAC5,
32'hBC8FEE89,
32'hBCD6F810,
32'h5CF1832,
32'h3D87FB13,
32'hBD10AA2C,
32'hBD08E90E,
32'hBD5B213A,
32'h3DB8B8EA,
32'hBDCAC8B0,
32'hBD627215,
32'h3D935CDC,
32'h3D7E44A1,
32'h3E00BC4C,
32'h0EC84BF6,
32'hBDD16142,
32'hBD184335,
32'hBDBE8648,
32'hBD07A41A,
32'h3EE5E369,
32'h3E8C39C0,
32'h3E1C707D,
32'h0EDEB349,
32'h3D7C42AB,
32'hBD38509D,
32'hBE9D9C0D,
32'hBE64062A,
32'h2ED2345F,
32'hBF0A83C2,
32'h3D440692,
32'h3CF18367,
32'hBEE9E04D,
32'h3DEEDF3B,
32'hBD6F4210,
32'h3E7F2D9F,
32'h3C2459B5,
32'hBF5038FB,
32'h3F5FBFC3,
32'hBE1C20A8,
32'h3F22BECE,
32'hBD3605BB,
32'h3EB65DDE,
32'hBCA87F35,
32'h3E13C0CA,
32'h3E9F51CA,
32'h3FA4735D,
32'hBEE10B24,
32'hBE610A9F,
32'hBE0751BA,
32'h3ED8D2B8,
32'h3EDA4772,
32'hBE3EC6E5,
32'hBC166D3F,
32'h3CA3261D,
32'h3D6242C0,
32'h3E3DA581,
32'hBE0F6F1F,
32'h3EC4E47B,
32'hBDA8757B,
32'hBEBE4E3A,
32'hBE147842,
32'hBF888917,
32'h3F63A635,
32'h3CD4FEE2,
32'hBE9063F7,
32'h3DC9385D,
32'hBF495277,
32'h3F613182,
32'h3EB87C3F,
32'h3DAE0F73,
32'h3EB09FEB,
32'hBF002222,
32'h3F9FB94F,
32'h3F170266,
32'h3EB57CED,
32'h3EBC57AE,
32'hBF896EB3,
32'h3EAD5F13,
32'hBE32E4BB,
32'hBE3EEB23,
32'h3EB4FF50,
32'h3F4F0FF9,
32'h3D21DD70,
32'hBE0CC67E,
32'hBD84E90C,
32'h3D0725B2,
32'h3C02F1ED,
32'h5DC851F5,
32'h3F003D72,
32'h3E2E87F9,
32'hBEB2E51B,
32'hBFB5192D,
32'h3E3E94EC,
32'hBEBF3A40,
32'h3E784C21,
32'hBE8E7A9D,
32'hBEE36DD9,
32'h3EEDC88F,
32'h3E9F1430,
32'h3EF1E5BE,
32'h3ED5FAD1,
32'h3DD07C48,
32'hBE8CD8AE,
32'h3EB1BE8A,
32'h3E917A0D,
32'hBFA5856E,
32'h3ECFDE06,
32'h3EEA0FB2,
32'h3DCF9AC1,
32'hBF2DD3CF,
32'h3E8FE459,
32'h3EB342D6,
32'hBC532C5A,
32'hBCE36887,
32'h3CF38CB4,
32'h3CAE9202,
32'h3E638781,
32'h3C8E1C01,
32'hBD092694,
32'h3DBC43EC,
32'h3E2179FE,
32'hBD0CF710,
32'h3E70E0EC,
32'h3EAB3BA7,
32'hBE9373C6,
32'hBF34A784,
32'h3D213C26,
32'h3CE8102B,
32'h3E348D61,
32'hBDB8C154,
32'h3E14CAB9,
32'h3DA72540,
32'hBEED1BE5,
32'hBEAC2162,
32'hBDA05E91,
32'hBF80D5F8,
32'h3D84A52F,
32'h3F17233E,
32'h3E85B927,
32'hBE975A32,
32'h3E518AF8,
32'h3E740DC3,
32'h3F82198A,
32'h3C83AA64,
32'h1DFD72D0,
32'h3C9181AC,
32'h3DFEBEA3,
32'h3DC84348,
32'h3E97C2F2,
32'hBD44A411,
32'hBE6558ED,
32'hBD99737F,
32'hBDA8989B,
32'hBEBE886A,
32'h3F0194AB,
32'hBE40F85B,
32'h3F1FF3E1,
32'h3DD86D68,
32'hBE69FE96,
32'h3E260CBB,
32'h3F43B9EF,
32'h3E59F8EF,
32'hBE7FFC7B,
32'hBEAC348B,
32'hBEDE8C54,
32'hBF8CB1B7,
32'h3E5C58C1,
32'h3E126D95,
32'h3E61FC62,
32'hBEABEDC3,
32'h3E7E3433,
32'h3F549849,
32'hBE83E889,
32'hBC580A72,
32'h3C111D05,
32'h3E1BF997,
32'h3F089205,
32'h3EB819DC,
32'h3EB3FEF6,
32'h3CDDB983,
32'hBD857C23,
32'h3C22B875,
32'h3DD36FC6,
32'h3DEB8B5A,
32'h3D6698AA,
32'hBF3665C8,
32'h3E10BD2D,
32'hBEB8840E,
32'hBF88EE0D,
32'h3DB3253B,
32'h3E36E23C,
32'h3E9BC256,
32'h3E65AC3F,
32'hBE32908A,
32'h3E5F070E,
32'hBF25E472,
32'h3EC105E5,
32'hBE43F2C1,
32'hBDBE53F0,
32'hBE6AD79F,
32'h3E347D2B,
32'hBE434CC1,
32'h3D3C7119,
32'h3D323884,
32'hBDB66F5F,
32'h3DB4D9EE,
32'hBE2CEBD1,
32'hBD3F3973,
32'h3E62CB9D,
32'hBEA22F7B,
32'h3E54BDFB,
32'h3EE1098E,
32'h3EB24664,
32'hBEA407A6,
32'h3E45EDBC,
32'h3D57200A,
32'h3E9679D5,
32'hBE8E00D3,
32'hBF782A63,
32'h1DECF1C5,
32'hBEADE234,
32'hBD6E3EC1,
32'h3EE2994A,
32'hBECBC645,
32'hBE8AE9C6,
32'h5DE0A8D7,
32'h3F083C64,
32'hBE667410,
32'hBF35B966,
32'h3DD32B9A,
32'h3DC416AE,
32'hBEE3E284,
32'hBDB7782F,
32'hBD724139,
32'hBC8ECF30,
32'h3D03165F,
32'h3E10A3D5,
32'h3EC03B85,
32'h3ED61C57,
32'hBDB2931A,
32'hBD844653,
32'h3ED8C355,
32'h3E8A1C08,
32'h3EB5569D,
32'h3D14D29A,
32'hBC8BFD6A,
32'h3ECF3856,
32'hBED9F721,
32'hBFB1825C,
32'h3C9231EB,
32'hBF10F729,
32'h3D9212CC,
32'h3E830D76,
32'hBE1B14C3,
32'hBE9B5987,
32'h3F089547,
32'h3F1D6048,
32'hBEB3C723,
32'hBF74D9FB,
32'hBF1EBCE5,
32'hBD2DCB34,
32'h3E1033EE,
32'h3E6C7651,
32'hBDC23971,
32'hBCDBF97D,
32'h3E0E102E,
32'h3E101739,
32'h3E34E5F3,
32'h3E93F481,
32'hBC35ED4C,
32'hBE444E55,
32'h3C6B207D,
32'h3E2387C3,
32'hBD8DC8AB,
32'h3CEDDB81,
32'h3DBDFD10,
32'h3E9A8056,
32'hBE08E818,
32'hBF27C2C3,
32'h3D8DB3F5,
32'hBE49FFEF,
32'h3E523F1E,
32'h3E74592B,
32'h3D15CA98,
32'hBDF9CC14,
32'h3EB029CB,
32'h3F275BA6,
32'h3E5D7CC0,
32'hBF696AE0,
32'hBF8801CC,
32'hBD416EDB,
32'h3E4ED806,
32'hBEAA12CC,
32'hBDC1CEDD,
32'hBDA8B56F,
32'h3E41FBF4,
32'h3E976668,
32'h3D887FB0,
32'h3EB422B5,
32'hBD6AB57F,
32'hBD93674F,
32'h3E90A411,
32'h3DA3A89A,
32'h3D6A82C1,
32'h3C5EE230,
32'h3EEB0442,
32'h3E25E6D5,
32'hBE30F21D,
32'h3EF9E60B,
32'hBD5BF79A,
32'h3E1B0FAD,
32'h3E249163,
32'h3F0FE52B,
32'h3E804B10,
32'hBFB068C9,
32'h3E85A80C,
32'hBE6C5F33,
32'hBDA95B53,
32'hBF6EEF41,
32'hBFBF2FF4,
32'hBEA37243,
32'h3E094160,
32'hBE92FD2D,
32'hBD9279E7,
32'h3C49126B,
32'h3E97BB8E,
32'h3DEC7ABB,
32'h3E0530E8,
32'h3C4A2ED2,
32'h3D1F8A49,
32'h1DEE2FA9,
32'hBC99CF09,
32'hBE9025D3,
32'hBEB64C19,
32'h3C856784,
32'h3E16EB6C,
32'h3DFD771D,
32'hBDE01EF8,
32'h3E1D3772,
32'h3E6D9B4F,
32'h3E724205,
32'h3DBB8F1A,
32'h3DF851A4,
32'h3ED6FEC0,
32'hBFF25634,
32'h3D9DC6D6,
32'hBF8A6494,
32'h3DE488A5,
32'hBECE1018,
32'hBFC771EB,
32'hBEF04107,
32'h3D5EEE3F,
32'hBDA87C19,
32'hBC330712,
32'hBD0BACB0,
32'h3E1C37BA,
32'h3E511EFC,
32'h3DCCEC4F,
32'h3E1E4C6F,
32'h3DF3AC71,
32'h3D077C43,
32'hBE75DBCA,
32'h3D1AACD9,
32'hBE827742,
32'h3D7AFCBB,
32'h3ED81C29,
32'h3E8E1A64,
32'h3E3DC41B,
32'hBE9C0D26,
32'h3F05E968,
32'h3DDAB2C7,
32'h3D2F5503,
32'hBEF27C60,
32'h3E135B71,
32'hBEF76D17,
32'h3E231636,
32'hBF5FBB7F,
32'h3E93286C,
32'hBEBB1F71,
32'hBF6E68C1,
32'hBEEFC171,
32'h3E02D47C,
32'h3EB24E41,
32'hBD9E67AF,
32'h3C909C1B,
32'hBC8899F8,
32'h3EA6189F,
32'hBE23AEB1,
32'h3EE437D3,
32'hBD3DA70C,
32'h3E2D57E4,
32'hBE6230EA,
32'h3E116368,
32'h3E0A001B,
32'h3E8D5B9A,
32'h3DD3A270,
32'hBE598F3B,
32'h3EA12B6F,
32'h3E045531,
32'h3E9BB9BE,
32'hBE306885,
32'h3E7D40E3,
32'h3E65D35B,
32'h3D8A4A05,
32'h3E9F7BA2,
32'h3EAC606F,
32'hBF5FF3FD,
32'h3C06EAF7,
32'h3D1B74C6,
32'hBF577783,
32'hBEED3393,
32'h3D898AB8,
32'h3F01039B,
32'h3CA8E9D1,
32'hBD709D33,
32'h3E3F2CAE,
32'h3EC8F063,
32'hBE80DBDC,
32'h3ED17A73,
32'hBD51FF46,
32'h3DAAD48E,
32'h3E03738F,
32'h3E355AB6,
32'h3D030CBC,
32'h3DD2EC43,
32'hBCFE9F4B,
32'hBD835536,
32'h3E5C78AC,
32'h3D84D7E0,
32'hBE113D81,
32'hBECD4734,
32'h3E1F461B,
32'h3E893702,
32'h3D9DCA76,
32'hBE71AB33,
32'h3DC01A94,
32'hBEE63283,
32'h3DA6AA4F,
32'hBE4D3478,
32'hBEADEC50,
32'hBE41D750,
32'h3DA6AB94,
32'h3E277372,
32'h3D21F307,
32'h3D08660D,
32'hBD8331F8,
32'h3D6814D9,
32'hBE3DC155,
32'h3ECA668C,
32'hBF25188B,
32'h3D994940,
32'h3E94FE3C,
32'h3D9FA3CF,
32'hBD368F3B,
32'h3E859F54,
32'h3E20AF5B,
32'h3C0CF53E,
32'h3E7726C8,
32'hBD3DA72A,
32'hBE923382,
32'h3CF04AB9,
32'h3DDAC89E,
32'h3ED8A177,
32'hBF09862A,
32'hBD61617D,
32'h1DFF0553,
32'hBD37FEBF,
32'hBC7CFF01,
32'hBE2342EA,
32'hBD073A80,
32'h3D382EC2,
32'hBDDD73AC,
32'hBD90C6D4,
32'h3CB93540,
32'hBD2C35BB,
32'h3E0AA126,
32'h3DD64E3C,
32'h3E0C8DD9,
32'h3E4CE2AF,
32'hBF8690EC,
32'h3E9DE4DB,
32'h3E209CBD,
32'h3E1222EF,
32'h3E86EE2C,
32'h3E2106BF,
32'h3E98C40B,
32'h3DAB3DD3,
32'h5DC4FED2,
32'h3E4AD3BE,
32'hBE9B74F6,
32'h1DF15E98,
32'h3DA0D006,
32'h3E7BE495,
32'hBED7A24E,
32'h3CAF9020,
32'hBE0BDB79,
32'hBD9B8B71,
32'h3DBBEE4D,
32'h3D5F1310,
32'h3DA3A55E,
32'h3DAD2B42,
32'hBCD637B9,
32'hBF46D6C5,
32'hBDD59E82,
32'hBD7F6E17,
32'h3ECBC436,
32'hBD4B255E,
32'h3DB9BDF1,
32'hBD37A612,
32'hC0050062,
32'h3CDBF64C,
32'hBC477994,
32'h3EFAB88E,
32'h3E05BA56,
32'h3ED18305,
32'hBD00F31F,
32'h3D62F446,
32'hBD090557,
32'hBE1E20DD,
32'hBE7D7BBE,
32'hBE1975F3,
32'h3D9F8091,
32'h3E20B813,
32'h3EEA99BF,
32'h3D3DFA8F,
32'h0EC5B2CF,
32'h3DA2DE87,
32'h3D4B57DE,
32'h3E9879F9,
32'h3E59AAE6,
32'hBE2E203F,
32'h3DE3B6D1,
32'hBED066C9,
32'h3CA219FE,
32'hBD58E77D,
32'h3EA9D610,
32'h3D225DD5,
32'h3D31B0F6,
32'hBDABBFD6,
32'hBFB3BBD7,
32'hBD15398E,
32'h3E3FB277,
32'h3E6A425E,
32'hBDD43FF4,
32'h3E904452,
32'h3D9F6289,
32'h1DFDA24B,
32'h3E01A401,
32'h3EC607FD,
32'hBE06EEE3,
32'h3E39D282,
32'h3E5BE662,
32'h3E12F3A6,
32'h3E62AAEB,
32'h3D961752,
32'hBDAC8A70,
32'h3DBF2FE4,
32'hBE1FCFF1,
32'h3DF61D64,
32'h3ECC3B0C,
32'h3DB39B54,
32'h3E91A212,
32'h3EB7591D,
32'h3C9B23BF,
32'hBDC0DD3F,
32'h3DB1D64E,
32'hBD578EE6,
32'hBE49D6DE,
32'hBD48ED01,
32'hBD274DA5,
32'h3E543545,
32'hBDE65D96,
32'h3EE0AC65,
32'h3D420A6F,
32'h3F00B110,
32'h3EA878AA,
32'h0ED114F9,
32'hBDD8BB9D,
32'hBD047A13,
32'h3C051C60,
32'hBDB6BD11,
32'h3E72BE14,
32'h3EFFB25C,
32'hBD95647C,
32'h3E22050E,
32'hBE6C9246,
32'h3EA17AD6,
32'h3C9CE52C,
32'h3E89180F,
32'h3E2882C7,
32'hBE317299,
32'h3E9D3055,
32'h3EB19602,
32'h3CD5C6A7,
32'h3C56890E,
32'h3E8D3BEC,
32'h3E0375CC,
32'hBDA6BDB4,
32'hBD59103C,
32'h3F091289,
32'hBEF2D041,
32'hBCABFE79,
32'h3F02DE2F,
32'h3F06E56D,
32'h3F1456CF,
32'h3E270FC2,
32'h3E3C494A,
32'h3D231D27,
32'hBE8CBF2D,
32'h3D2E2CE6,
32'h3CCFE9D6,
32'hBD2D4C7A,
32'h3F066530,
32'hBDEB66B3,
32'h3EAC2DC5,
32'hBE876B29,
32'hBD43F0DE,
32'h3E9A9B04,
32'h3D369283,
32'h3EB3EBF3,
32'h3EEB912C,
32'hBD6F501D,
32'h075FF4B0,
32'h3D4311E0,
32'h3D1FED36,
32'h3E0FEE00,
32'hBE9DD054,
32'h3EA38706,
32'hBE13D997,
32'h3EEDAD56,
32'h3E4286A1,
32'hBE5CEA55,
32'h3E64D06C,
32'h3EF11439,
32'h3EA37B66,
32'h3E47AA81,
32'h3D89C57A,
32'hBD99F5EA,
32'h3DE53B57,
32'h1751C523,
32'hBEEAC3C2,
32'h3CA20066,
32'h3F128DB8,
32'h3DF3EB8E,
32'h3E7D9A1C,
32'hBEA30889,
32'h3D704A88,
32'h3E2C4080,
32'h5DE92795,
32'h3E8C274D,
32'h3E0DC756,
32'hBEDB88FE,
32'hBE7B9DBA,
32'h3D1D8607,
32'hBC3F5A67,
32'h3EEC2F1A,
32'h0ECA4476,
32'h3E157690,
32'hBD80BF3C,
32'h3E519B74,
32'hBE84670D,
32'hBE10840B,
32'hBDC44C93,
32'h3F18BC0F,
32'h3E07A788,
32'h3DAF8074,
32'hBE257C54,
32'hBEC31566,
32'hBE950EEA,
32'h3DCB6F7C,
32'hBF90E34D,
32'h3DF5E08B,
32'h3EB8B30C,
32'hBD3ECF89,
32'h3C08C6A3,
32'hBE5CDDA1,
32'h3D597071,
32'h3DBDF9CB,
32'hBDD6C2BC,
32'h3EA40D07,
32'hBE4F3420,
32'h3D219B20,
32'hBE3F6904,
32'hBCFA84DB,
32'hBDEBCA89,
32'h3E684111,
32'h3E5B9E5D,
32'h3D0733DB,
32'h3D9C99D2,
32'h3EAE0135,
32'hBEF879EC,
32'hBE88A7A6,
32'h3EDC1A04,
32'h3F14FF68,
32'h3DC7AF72,
32'hBF263A93,
32'hBE59E131,
32'hBEE8BECE,
32'hBEC5818D,
32'hBE703DF5,
32'hBF8DD4D4,
32'h3EDF2A94,
32'h3ECA5DED,
32'h3F284FE8,
32'hBEA2F89A,
32'h3EBB6D5B,
32'hBE11EDC9,
32'h3E0B2AA7,
32'h3F153130,
32'h3E12EFE0,
32'hBE5D1FCB,
32'h3DA5230E,
32'hBF006220,
32'h3C757C79,
32'h3CD9F81C,
32'h3DC7BB78,
32'h3DE321A8,
32'hBEB3DE1C,
32'h3DC63533,
32'hBEEC53DA,
32'hBE8F50A8,
32'hBEED34D0,
32'h3E6D1AA4,
32'h3EE5475C,
32'h3E5B0898,
32'h3E4B01DF,
32'h1DDBBFD2,
32'h3E401FCE,
32'h3D899694,
32'h3EFE5AC2,
32'hBEFA2B4B,
32'h3E76D32F,
32'h3F307874,
32'h3F31A218,
32'hBF0A9F28,
32'h3F5D6F61,
32'hBF14BE88,
32'h3F5A4970,
32'hBFA7C078,
32'h3ECED376,
32'h3F01EE22,
32'h3F295BF9,
32'hBC9E8CD6,
32'hBDBB9344,
32'h3C172E8E,
32'h3F3D8A0D,
32'h3F1E0F57,
32'h3FAB0B58,
32'hBDD9C10E,
32'h3EC09DCD,
32'h3F015A63,
32'hBF8D5394,
32'h3F423B59,
32'h3F671E1A,
32'hBED2FA61,
32'hBF18331F,
32'h3DCC666A,
32'h3F6AD1EB,
32'h3EA3A926,
32'h3D8661F5,
32'hBF28C532,
32'h3F38E225,
32'hBE43616F,
32'h3E9E739A,
32'hBE1EE9F9,
32'h3F594722,
32'hBFBD2CFC,
32'h3F0CAF05,
32'hBF8F6C88,
32'h3EDE3F84,
32'h3DFCA5FB,
32'h3F3BBC12,
32'h3EA6D321,
32'hBDA50C0A,
32'h3CCDF597,
32'hBEA2B183,
32'h3F90E3A6,
32'h3F76ADE7,
32'hBE92DA6E,
32'h3FA5A850,
32'h3E03219C,
32'hBFAF918B,
32'h3F46C28C,
32'h3F10B902,
32'hBF03E80E,
32'hBF78AA7C,
32'h3E0E343D,
32'h3F245B0A,
32'h3E0264FE,
32'hBE395314,
32'hBEF2751F,
32'h3F012B57,
32'hBF02C0ED,
32'h3CA5B6BF,
32'h3D040451,
32'h3F31AEEE,
32'hBF5C4301,
32'hBDF29747,
32'hBE32885E,
32'h3FC81395,
32'h3F240425,
32'h3F82387D,
32'h3F05F223,
32'hBD8E032D,
32'h1DCFE2CE,
32'hBDA2859A,
32'h3F97F57C,
32'h3E1D6407,
32'hBF45102E,
32'h3FC4157F,
32'h0EC61966,
32'hBEEA851D,
32'hBF1BDBDB,
32'hBE490B04,
32'hBEC7D875,
32'h3DF1CB35,
32'hBF81630D,
32'h3F860119,
32'hBCD411FE,
32'h3FC7A06C,
32'hBEDD6C45,
32'h3F140224,
32'hBF967308,
32'hBD7D96CE,
32'h3F1F2700,
32'h3D02055E,
32'h3CFE472F,
32'h3D992867,
32'h5DC4FB1D,
32'h3F5636D5,
32'h3ECE8251,
32'hBC8F07CD,
32'h3D22CEEF,
32'hBD3BE8CA,
32'hBCDD50DD,
32'hBD9C45E9,
32'hBD8F7DB9,
32'hBCDFA5F2,
32'hBF0D537D,
32'h3DBB6CC9,
32'hBE17FD6E,
32'h3F4DA09B,
32'hBC112FE1,
32'hBF9A8749,
32'h3F187460,
32'h5DE17709,
32'hBF8123E2,
32'hBD93C323,
32'h3EB46F78,
32'h3F4BEE2C,
32'h3ECCFA26,
32'hBCF167A1,
32'hBF6A820F,
32'h3D0204D5,
32'hBC9FAD84,
32'hBDB026A0,
32'h07594F88,
32'hBD90BF5A,
32'hBDB8162C,
32'h3F0C15ED,
32'hBE5B0942,
32'h1DC59210,
32'h3D183C18,
32'hBC9E7671,
32'hBD89DDBE,
32'hBE6CE88D,
32'hBD986F35,
32'h3C9076B7,
32'hBEA1C2E4,
32'h3E0743C7,
32'hBD86DD1C,
32'hBE732BF7,
32'h3D7C84AB,
32'h3D9F156C,
32'h3CBB8EE7,
32'h3C320E0F,
32'hBEE52689,
32'h3EDB4670,
32'hBD9B9095,
32'h3DDD57D4,
32'hBD9D8F23,
32'h3E28E85F,
32'h3D2B0174,
32'h3D36E376,
32'h3EC591E8,
32'hBCF1CF85,
32'hBF318B1A,
32'hBEA6C89F,
32'hBED57350,
32'hBD75F13A,
32'hBEC49F27,
32'hBEED9F32,
32'hBDB8413B,
32'hBDCE7D4D,
32'h3D801C43,
32'h3DC41BDB,
32'hBF09CC08,
32'h5DC61C2D,
32'hBD8C91E7,
32'hBEA32284,
32'h3D8561AA,
32'hBF580F33,
32'h3F36BA8A,
32'h2ECB38AC,
32'hBE102D14,
32'hBD60617E,
32'hBED1C763,
32'h3E99935D,
32'h3ED8260C,
32'hBE797680,
32'h3E0CD048,
32'hBF3DCD23,
32'h3FBFAC0D,
32'h3F1CF34D,
32'hBEA0F00C,
32'hBF1E75D3,
32'hBF9441AF,
32'h3EAB3B7B,
32'hBF0C3577,
32'h3EFD7277,
32'h3EF88EFA,
32'h3E263625,
32'hBE9F6F07,
32'h3D16EDC4,
32'h3D708BB6,
32'hBF13E4BE,
32'hBE43CB7A,
32'h3E8DF4D3,
32'h3E1557FC,
32'hBDA4BDCC,
32'h3F1E79C5,
32'hC011FC51,
32'h3E905D52,
32'h3F6B7CC0,
32'h3DE89301,
32'hBF04364F,
32'hBF1C5902,
32'h3F57766A,
32'hBF83C09C,
32'h3ED69FE6,
32'h3EA454D7,
32'h3E4D97F8,
32'h3F049D56,
32'hBEAEC996,
32'h3EFF89B0,
32'hBF023621,
32'h3C9444C2,
32'h3E954296,
32'h3F057619,
32'hBF455E3F,
32'hBDF7E5C3,
32'h3E8A0EFC,
32'hBDEBBA75,
32'hBD0D158E,
32'h3D46F9EC,
32'h3ECD231C,
32'hBE06A15C,
32'hBCFEFE55,
32'hBC9D3B21,
32'h3EEB896B,
32'h3E54F2FD,
32'hBF21672E,
32'hBD504EA1,
32'h3F0C9396,
32'h3D9F40B6,
32'hBF245C7A,
32'h3EBB9E5F,
32'h3EAB95DE,
32'hBE431616,
32'h3EDCA900,
32'h3E526F5A,
32'h3EC836D2,
32'h3E82B3EA,
32'hBF93A2D4,
32'h3EA30732,
32'hBED93C1D,
32'h3E293439,
32'hBCEAEA21,
32'h3E9AF3EE,
32'h3E780B92,
32'h3F079C12,
32'h3E8182D0,
32'h3D983B1A,
32'hBC854086,
32'h3DAA5A9F,
32'hBE209B0E,
32'hBD809648,
32'hBC8CB9CC,
32'h3DBFA617,
32'hBF4322E6,
32'h3D0C62E2,
32'h3DCFFD01,
32'h3DC0DC46,
32'hBE47DC8F,
32'h3E84082C,
32'hBEFA52CE,
32'h3E9EA256,
32'h3C778477,
32'hBE0F07AB,
32'h3E80C356,
32'h3E5D0ED5,
32'h3ED5286B,
32'hBE9F0A9E,
32'hBF4B3BB0,
32'h3E4FB38F,
32'hBE25C9FF,
32'h3E355414,
32'hBDFE230C,
32'h3E3ECA75,
32'h3F0F97FC,
32'h3E9B57B9,
32'h3E96FEB6,
32'hBFACAA68,
32'hBCA4293A,
32'h3C9351C3,
32'hBD1A4675,
32'h3F05EA5D,
32'h3E232518,
32'h3E0BD7E0,
32'hBEBD746F,
32'h3E561418,
32'h3E30BFC4,
32'h3E91EE31,
32'hBCCB105E,
32'h3E9AD3EE,
32'hBFA175AB,
32'h3E476AB4,
32'hBEA48EC2,
32'hBED81CD1,
32'h3C62F73D,
32'hBDAB0B1E,
32'h3DB9A13B,
32'h3D9C7B7F,
32'hBEEFEE3F,
32'h3E9A1E79,
32'h3F04377F,
32'h3E9448F0,
32'h3DC96E1C,
32'h3EEDDD9C,
32'h3E83BC16,
32'h3E9078FE,
32'h3D740D34,
32'hBEA59FD0,
32'h3CC10C39,
32'h3D1186A4,
32'h3EAC726F,
32'h3ECF1B07,
32'h3E3F700B,
32'h3E326564,
32'hBE953204,
32'h3E51EF29,
32'h3F0C95E1,
32'h3ED00712,
32'hBEAE8467,
32'hBE14FC70,
32'hBE715199,
32'h3EE65819,
32'hBEF81065,
32'h3D69A809,
32'hBEB1C863,
32'hBEE08866,
32'h3E1DA564,
32'h3F062C7A,
32'hBDFADFE7,
32'h3EC59BD7,
32'hBE5F22FB,
32'h3F0E1893,
32'hBE866468,
32'h3EE3BB11,
32'h3E445D37,
32'h3F025B5D,
32'h3D664FC9,
32'h3DDE410C,
32'hBD4E5507,
32'h3C518A20,
32'h3E0B782E,
32'h3EC60840,
32'h3EBFACD2,
32'h3E82C295,
32'h3E29910D,
32'hBD601C9E,
32'h3E40CA68,
32'h3E9C1587,
32'hBF104970,
32'hBC8C1D32,
32'hBD8A3F32,
32'h3F09812B,
32'hBF075A62,
32'hBE4BD9CB,
32'hBE27C90C,
32'hBF1B21E9,
32'h3E8E805A,
32'h3D823EB1,
32'h3D0DE832,
32'hBE4C1338,
32'h3D4C1D76,
32'h3F2A7EB1,
32'hBF1A8B7A,
32'hBE7F1465,
32'h3D092A60,
32'h3F128BD3,
32'hBCC64052,
32'h3DA6E9A2,
32'h3C4DF9F7,
32'h3D1C0668,
32'h3DEF3B23,
32'h3E513881,
32'h3E972C92,
32'h3F330B3C,
32'h3EA9D822,
32'h3E459619,
32'h3EA6CAD6,
32'h3E9FB153,
32'hBF08250A,
32'h3E316E8A,
32'h2EC728B2,
32'h3EF32917,
32'hBCE8831C,
32'h3E4B83AC,
32'hBE240BA4,
32'hBF14151C,
32'h3D8351CD,
32'h3E96CB3B,
32'h3E21DF82,
32'hBF6C8A7E,
32'h3E38ED46,
32'h3F137378,
32'hBE26C0E2,
32'hBF1C3549,
32'hBE1B09AC,
32'h3EF67E63,
32'hBE1FE697,
32'hBDAE3EC0,
32'hBC63866A,
32'h3CD2132B,
32'h3ED0304E,
32'h3D05B4BD,
32'h3E0FF964,
32'h3F5A0E8A,
32'h3EB02555,
32'hBD6BB8F3,
32'h3EC1D734,
32'hBE3BDF3E,
32'hBE541E96,
32'h3E9BE71A,
32'h3E55A3C0,
32'h3F019A2E,
32'hBEF6CB45,
32'h3ED94738,
32'hBDDB8756,
32'hBEC85AD6,
32'hBE20C4F0,
32'h3EFDFEE6,
32'h3EC5B1ED,
32'hBFA7A046,
32'h3ED35510,
32'hBD34E22E,
32'hBE898798,
32'hBF059363,
32'h3C26B75C,
32'h3EFF20F3,
32'hBD7C51D7,
32'hBE4C4ACC,
32'hBD7AB29E,
32'hBDB1165D,
32'h3EAF5E4C,
32'h3E826E26,
32'h3E58F204,
32'h3F57A35E,
32'h3F137AF8,
32'hBE1CC4CC,
32'h3DD8D20A,
32'hBE8C6EED,
32'hBC2FA5C5,
32'h3E6849DF,
32'h3ED2FEA8,
32'h3F2B25BD,
32'hBED078C9,
32'hBE0235F4,
32'h3DC191E4,
32'hBE6F36CB,
32'hBE4F8E18,
32'h3E08DBBA,
32'h3EC7F044,
32'hBF03EC54,
32'h3EA6C184,
32'hBF4F5C3F,
32'h3E8CBD6D,
32'hBF345E61,
32'hBE706091,
32'h3F34140A,
32'hBC82B9CC,
32'hBE843BFD,
32'hBC3FA13D,
32'h5DF0A59B,
32'hBD7FC645,
32'h3E8B990A,
32'h3E854174,
32'h3F494FEB,
32'h3E5D5A87,
32'hBD8AFD22,
32'hBE2D91C9,
32'hBE096205,
32'h3DB701F6,
32'h3EBB8ADB,
32'h3F10F07D,
32'h3F2984FD,
32'hBDC272BA,
32'hBE894105,
32'h3E3F2F4F,
32'h3E6D9866,
32'hBE0B456A,
32'h3EEE3DAC,
32'h3E6E9855,
32'h3EDB0175,
32'h3EC6A550,
32'hBF1219E0,
32'h3EB20F91,
32'hBE253DFD,
32'hBF197158,
32'h3ED91913,
32'hBE9925F0,
32'h3E92F0A0,
32'hBD720053,
32'hBD9565EB,
32'h3E7FC8B4,
32'h3E9E50D9,
32'hBC3A3C5F,
32'h3F28A5C9,
32'hBE577843,
32'h3E82D12A,
32'h3E84A709,
32'h3E02E28B,
32'h3D691537,
32'h3E90D0A5,
32'hBE9BF6A1,
32'h3E860FBC,
32'hBE164D7A,
32'h3EAF6EF2,
32'h3D027F5B,
32'h3D63A70F,
32'hBDA666B3,
32'h3F225597,
32'h3C008657,
32'h3EF06E96,
32'h3E9DB76B,
32'hBEC7D2D0,
32'hBE16B144,
32'hBCE04858,
32'hBF1D298E,
32'h3E2DA3BB,
32'hBD96D005,
32'h3EE06B16,
32'hBE37B7D1,
32'h3CE5B5F1,
32'h3EFAD60C,
32'h3E78CC8D,
32'h3D5F0C3A,
32'h3E9D465E,
32'h3D154B1B,
32'h3E17343C,
32'h3EAF9105,
32'h3D83CDB7,
32'hBE489CB8,
32'h3DB2E7D9,
32'h3E9CD24A,
32'h3EE8FA64,
32'hBDB07292,
32'h3EDA1B14,
32'hBEB41AAA,
32'hBDD7B8B1,
32'hBD8413C4,
32'h3E2137EE,
32'hBEE6376B,
32'hBE12FD75,
32'h3E1EB43B,
32'h1DDDFE0B,
32'hBDD046AF,
32'h3D66EF23,
32'hBE3AF730,
32'h3D3578C5,
32'h3C798EA9,
32'h3D62D2EE,
32'hBDF8A6C0,
32'hBD850547,
32'h3E59FE75,
32'h3DC339EE,
32'hBC0CAB61,
32'h3EB66B7F,
32'hBF80943F,
32'h3C98767E,
32'h3E1FE8B6,
32'hBCFEF9C5,
32'hBD01215F,
32'h3E6BD223,
32'h3EA81A01,
32'h3EA9A939,
32'h3E0D3798,
32'hBE671D08,
32'hBE72CD38,
32'h5DD38D99,
32'hBD90224C,
32'h3DFAD618,
32'hBF3060AB,
32'h1DF978A5,
32'h3E0488AF,
32'hBCFBD331,
32'h3E7378C1,
32'h3DC080CA,
32'h3E280A00,
32'h3CC5433B,
32'hBE62269E,
32'hBEBB61B4,
32'hBD9F9406,
32'hBD871D70,
32'h3E1DE0B8,
32'h3E4BDB17,
32'hBD5AD649,
32'h3D1CA9CE,
32'hBF8F7823,
32'hBE23750A,
32'h3D7DFE33,
32'h3E14512C,
32'hBE4C5A02,
32'h3E918248,
32'h3EC3CB4B,
32'hBC358171,
32'h3E66FDFE,
32'h1CE89BA,
32'hBDFDC8EF,
32'h3E013718,
32'hBD41FBDA,
32'hBCB01573,
32'hBF0236F5,
32'h3D2F7EE3,
32'h3D819643,
32'h3E39629C,
32'hBE73BE52,
32'h3DDE3957,
32'h3E577127,
32'hBE03AD20,
32'hBD16B823,
32'hBE235637,
32'hBC27DCA6,
32'hBD5DDDCF,
32'h3EDF6728,
32'h2EDBE79F,
32'hBDE83920,
32'hBC70B75F,
32'hBF5731C0,
32'hBDDC64A5,
32'h3E03C852,
32'h3E0E5FFA,
32'hBF0C27A2,
32'h3DE9C780,
32'hBE7DF3D3,
32'h3E2CBE84,
32'h3E8D5158,
32'hBD99C32F,
32'hBE30756E,
32'h3EE356BA,
32'hBDA8ADD2,
32'h3DBC300D,
32'h3EAB75CC,
32'h3E5A9CD0,
32'h3E0732EE,
32'h3E424479,
32'hBE46C9B5,
32'hBDFB6F53,
32'h3E359470,
32'hBE8EE803,
32'hBD88D2C3,
32'h3E8A02E9,
32'h5DD9B184,
32'hBCF68A83,
32'h3E7F8051,
32'h3DF6E865,
32'h3E3DDFD7,
32'hBC7CB6D2,
32'h3DA9D212,
32'h3E01E84D,
32'h3D083002,
32'h3E8C132B,
32'hBE4AEC38,
32'h3DE2E31A,
32'h3CB8AEFE,
32'h3EA16B43,
32'h3E2A1EDF,
32'hBD89A2B1,
32'h3D742322,
32'h3EA04B82,
32'h3D794041,
32'h3E43D24A,
32'hBC38DB86,
32'hBC6902E9,
32'h3E45EDE7,
32'h3E080501,
32'hBEBED063,
32'hBDF23850,
32'h3EBD917A,
32'hBE319F38,
32'h3DB4CB99,
32'hBD8D7879,
32'h3D227B1F,
32'hBD3EA9F2,
32'hBDE71D6E,
32'h3DF1FF0B,
32'hBE2152F6,
32'hBD8D777A,
32'h3F17E9A0,
32'h3D12EB72,
32'hBDE4169B,
32'h3DFEBEF1,
32'hBF0882E0,
32'h3EB7081B,
32'h3EE86ACA,
32'h3E9F167D,
32'h3E7DF158,
32'hBECA076E,
32'h3E1D7D2E,
32'hBE5EB4D2,
32'h3E334AB8,
32'h3E89D70A,
32'hBFCA2188,
32'h3ECEE770,
32'h3CB09AD5,
32'h3DBAC39C,
32'hBEB8ED13,
32'h3D89EC52,
32'h3E9D7FDA,
32'hBE1CD4FA,
32'hBE28F657,
32'h3EBC2CCA,
32'hBD0D04F2,
32'h3C3F6996,
32'hBDB143EA,
32'hBE250BB0,
32'hBE85033A,
32'hBD7606A8,
32'h3EE74E71,
32'hBD3DEB60,
32'h0E496DE,
32'h3D5B79C3,
32'hBEF27A9F,
32'h3EC89424,
32'h3E491CE3,
32'h3D8F1B18,
32'hBD92E263,
32'h3E7AA63C,
32'h3E9B32EF,
32'hBCAE2553,
32'hBE39DF42,
32'h3DAE324B,
32'hBE586810,
32'h3F294852,
32'h3E540A7B,
32'h3E37F6EA,
32'h3E54751E,
32'h3E051DA5,
32'h3F7180F1,
32'hBE9A7949,
32'h3DB16669,
32'h3E824813,
32'h3C4D42DC,
32'h3C0FF2B1,
32'hBD2D3A08,
32'hBD8E7480,
32'h3E4C165B,
32'hBDD6A8D7,
32'h3F1FC632,
32'hBD1F574D,
32'h3DEA89B1,
32'h3E9C7141,
32'hBEB4E72C,
32'h3E2EB38F,
32'h3E3E338D,
32'hBDB24ED3,
32'h3D9C08E2,
32'hBEA74919,
32'h3DC1B36D,
32'hBE868675,
32'h5CC3E3F,
32'h3E868796,
32'hBF56F0AA,
32'h3F0F72E5,
32'h3D762443,
32'h3E4265B7,
32'h3DC4D30C,
32'h3D944053,
32'h3EFD2F7D,
32'hBE97611E,
32'h3E228370,
32'h3EAB1ED3,
32'hBD36A9A3,
32'h3CA8170A,
32'hBE301C6A,
32'hBD341202,
32'h3D9DAF74,
32'h3DCDD782,
32'h3F35BECA,
32'hBF09692B,
32'hBEFCE3BA,
32'hBE5EEA1D,
32'hBE406BB7,
32'h3E738BC1,
32'hBF500703,
32'h3D462ABB,
32'h0EC7937B,
32'hBF800F03,
32'h3E5E02CB,
32'hBE6E5DC4,
32'h3E1512EF,
32'h3E8D715D,
32'hBD9DCD62,
32'hBF2B09A8,
32'h3DA3D8F0,
32'h3DEE7B11,
32'hBE7F0798,
32'h3F11B50B,
32'h3D3B7065,
32'hBF3751EE,
32'h3E04A8DA,
32'h3EB690D0,
32'h3DDDEDAD,
32'h3DBBC382,
32'h3F16C496,
32'hBD732085,
32'h3D5D3DA3,
32'hBE1633B1,
32'h3F03AD02,
32'h3E5CDD95,
32'hBF760952,
32'h3E084D86,
32'h3E9425F4,
32'h3E9118E9,
32'hBF67F321,
32'h3E8BFFCF,
32'hBF0C0B3C,
32'hBF188D45,
32'h3DDD05D2,
32'hBF3595FB,
32'h3E54FF6E,
32'h3EC2D190,
32'h3E645FC0,
32'hBEF50DC1,
32'h3EE33FB5,
32'hBDC336CF,
32'hBEDAE829,
32'hBDCF3200,
32'h3C879C0F,
32'h3F1E9987,
32'h3EDEC859,
32'hBE272C68,
32'hBD450A46,
32'h3D98D3BD,
32'h3E6E67EC,
32'hBC99BA9C,
32'h3E2FEB76,
32'hBE784EAA,
32'h3E3C14B2,
32'h3DEE5AA6,
32'hBFA4A8C2,
32'hBDE4CDE5,
32'h3E934F1E,
32'h3EE72953,
32'hBFB503FE,
32'h3E6D7763,
32'h3E237314,
32'hBF16686F,
32'h3E8F5CAD,
32'hBEAD321C,
32'h3F00ABDC,
32'h3F23F581,
32'h3F2C8E05,
32'h3C248B52,
32'h3FA1AE53,
32'hBF3A4913,
32'h3EB6390C,
32'h3F223319,
32'h3EFA72E6,
32'h3F397751,
32'h3F857788,
32'h3F334427,
32'hBD101409,
32'h3CD595EE,
32'h3EE820B7,
32'h3F6F215E,
32'h3FA21D15,
32'hBDEB53BC,
32'h3F55358A,
32'h3E59C8D3,
32'h3DBDD987,
32'h3E4CD18C,
32'h3F03D074,
32'hBFA573D3,
32'hBFBF92C0,
32'hBF564D6B,
32'h3F93F981,
32'h3E90E01B,
32'hBF029D3B,
32'hBF03E7DE,
32'h3F2F46A6,
32'h3DF63CC9,
32'h3F124BE5,
32'h5CFC6DC,
32'h3F7560B2,
32'hBF7BDB03,
32'h3F68F935,
32'hBD895346,
32'h3E8A842B,
32'h3E134C34,
32'h3F3EEBF2,
32'hBDA997E8,
32'hBDB2ADCC,
32'h3E24A816,
32'hBF9E7517,
32'h3F82850E,
32'h3EBCFD7E,
32'h3E95CBDD,
32'h3FA8EABB,
32'hBCC29409,
32'h3DF0776C,
32'h3F1C3D12,
32'h3F97E113,
32'hBE2A2596,
32'hBEA14494,
32'hBF1AD72C,
32'h3F7C1A80,
32'h3E61BF92,
32'hBD7EF2A0,
32'hBE011A29,
32'h3F0A5B33,
32'hBED7AEAB,
32'h3F5EBCE5,
32'h3DD55318,
32'h3E1CBCF6,
32'hBF197C3B,
32'hBD60430A,
32'h3EDCEBD5,
32'h3F7C454A,
32'hBE332274,
32'h3F0A37C1,
32'h3FA90C03,
32'hBD3FD567,
32'hBD6A6F01,
32'hBECF2573,
32'h3F8210DA,
32'h3E161A50,
32'hBF4EEA06,
32'h3F6801C3,
32'h3D7AB3F5,
32'hBE97A7CE,
32'hBE6E750E,
32'hBEE90816,
32'hBF05ECCC,
32'hBEF3DD99,
32'hBFA24F76,
32'h3E925F55,
32'hBDFBBDC0,
32'h3F201FFC,
32'hBE3EBCA5,
32'h3EAA7106,
32'hBF17296A,
32'h3CF1F271,
32'h0EDAB88C,
32'hBD3DCC01,
32'h3D6B0372,
32'hBDA03C4A,
32'hBCB7E69C,
32'h3CD3F581,
32'hBD656783,
32'h3C7814BB,
32'h3D88B660,
32'h5DC109F9,
32'hBDDD0631,
32'h3D5A02F1,
32'hBC3496E7,
32'h3D0501A4,
32'h3C94FEC2,
32'h3E24B22A,
32'hBD2E1250,
32'hBD19B5E9,
32'hBCA16700,
32'hBDAFBE4D,
32'hBE15CCCC,
32'h3D1B36D8,
32'hBDFB1C35,
32'hBC7290DB,
32'hBD80F656,
32'hBD807B92,
32'hBDE3D454,
32'hBDB06303,
32'hBCA207DC,
32'hBD4CB53B,
32'h3F576999,
32'h3E2C1EE2,
32'h3D9FC5C7,
32'hBD108D5A,
32'hBDC29D7A,
32'hBC1049EA,
32'hBCBAD0E4,
32'hBC782CF8,
32'h3E1ED28C,
32'hBDBCA7FB,
32'hBD479CBD,
32'hBD72EC95,
32'hBE3F3CF8,
32'h3DE8D62D,
32'hBF43BDB4,
32'hBD228984,
32'hBC428A49,
32'hBD696F55,
32'h3D4C0F24,
32'hBF546FDC,
32'h3F930298,
32'h3C082776,
32'hBE238A83,
32'hBEFFFD41,
32'h3E8F5BE4,
32'h3EABDA28,
32'h3DA8EEE6,
32'hBD6B18E6,
32'hBF717E72,
32'h3F0010B9,
32'h3F4CE408,
32'hBDD09819,
32'h3FC6BF02,
32'hBECE99AC,
32'h3F915D32,
32'hBFAF7CC0,
32'hBEEAC757,
32'hBF1C6713,
32'hBDD134F3,
32'hBCECC051,
32'hBC8C31A5,
32'hBDF9B50C,
32'hBEF45176,
32'hBF137EDC,
32'h3E9574A0,
32'hBF178F18,
32'hBE8BAD3C,
32'h3EFD7200,
32'h3F1A291F,
32'hBF236A0D,
32'h3F1C3395,
32'hBE0485C8,
32'hBEBD596F,
32'hBEEC3DFE,
32'h3F7691A8,
32'h3FAC5DC9,
32'h3EE0E1B7,
32'h3E8A1C1E,
32'h3E81C9D4,
32'h3ECC1AFA,
32'hBF34B2CC,
32'hBF4EFB01,
32'hBEB41771,
32'h3EEC3AA9,
32'hBF33AD5F,
32'h3EB34C53,
32'h3F520134,
32'hBE3CB16A,
32'hBEB894C6,
32'h2EDF0873,
32'h5DDD81C5,
32'hBF1B07F3,
32'hBF517114,
32'hBDAC5810,
32'h3E2AE4F7,
32'h3F276B9B,
32'h3F5E22BD,
32'hBFD275D1,
32'h3EC134AB,
32'h3F5FC457,
32'h3EBBBF86,
32'hBED481EA,
32'hBD906746,
32'h3F057D52,
32'hBEDC59F6,
32'h3E3EF143,
32'h3E16D10E,
32'h3D7104BD,
32'h3F4E8C99,
32'h3D25997F,
32'hBD8A716C,
32'hBDC13C0E,
32'hBD298712,
32'h3DA6AAD9,
32'hBE7414B2,
32'hBE8486E1,
32'h3C8C7777,
32'h3EC826DA,
32'hBDACC70A,
32'h3D3E654D,
32'h3DA152CE,
32'h3E7E5744,
32'hBE413C63,
32'hBE0801C1,
32'hBD8CE848,
32'h3F3A7AED,
32'h3D77F679,
32'hBFFC2F18,
32'hBDAC77F2,
32'h3F5EBF1B,
32'hBD425B9C,
32'hBF58E3C2,
32'h3E439552,
32'h3E75B375,
32'hBE8B5B0E,
32'h3E0BC8A1,
32'h3F083195,
32'hBD88BC57,
32'h3E0D7C23,
32'hBF81B3E8,
32'hBE52EC26,
32'hBEB859C1,
32'h3EBCFDB1,
32'h3DB23308,
32'h3E2225C0,
32'h3EAD712B,
32'hBDB303A1,
32'h3EB785B5,
32'hBE4DEFCF,
32'hBD8A4401,
32'hBDB30AE2,
32'hBCCBAB5A,
32'h3D2AE244,
32'hBDCD63B7,
32'hBE9DD400,
32'h3DF44386,
32'hBCD5792E,
32'hBF382EFC,
32'h3E186DE0,
32'hBE4E5C10,
32'hBDC9C5B5,
32'hBFA668D6,
32'h3C8D7EEA,
32'h3E95E8FF,
32'hBCABFC01,
32'h3CA6D192,
32'h3EDA56DF,
32'h3E68C5D1,
32'hBED6A3AB,
32'hBF05F1B7,
32'hBE67CEC5,
32'hBDB88E80,
32'h3E1510A1,
32'hBEFF10CF,
32'h3E37D096,
32'h2EC92428,
32'hBE0860A8,
32'hBD3F8CE7,
32'hBFA4A71E,
32'h3C43610B,
32'h3D1C0B59,
32'hBCBAD8D7,
32'h3D6CE297,
32'h3EC61417,
32'h3D20B229,
32'hBEE4FE4B,
32'h3E28F786,
32'hBE2D07CE,
32'h3ECDEB95,
32'hBEDF4ED1,
32'h3E9FA9D8,
32'h3DCCEC01,
32'h3E157481,
32'hBDE57B7A,
32'hBF2F8A2B,
32'h3E3256E2,
32'h3ED558CC,
32'hBDF6EB08,
32'hBEA6F8FB,
32'h3E4A3348,
32'hBD3B40DF,
32'h3E6E1920,
32'h3E85EDCB,
32'hBE964753,
32'h3DAA248E,
32'h3E84C534,
32'hBD06D766,
32'h3D923CC8,
32'hBEA21FFC,
32'hBC9A2544,
32'hBD5F45FB,
32'h3E068058,
32'h3E73A877,
32'h3F1CC023,
32'h3E646FB5,
32'hBDCDDBC5,
32'hBEA048E2,
32'h3EB498FE,
32'h3E502074,
32'hBFBF1927,
32'h3DCD33B3,
32'h3E175F91,
32'h3E45B53C,
32'hBEBE4D58,
32'h3E0B07DA,
32'hBCECD74F,
32'h3E5F352D,
32'hBD73930C,
32'h3C8059E2,
32'h3DA71C97,
32'hBF07BF47,
32'h3C7A8F21,
32'h3E8BDD56,
32'hBEC0D51A,
32'h3E7B5593,
32'h3E5D669C,
32'h3DD985D2,
32'hBD8B9CCA,
32'hBF069402,
32'h3C654331,
32'hBCAE36E2,
32'h3E887D67,
32'h3E1BE742,
32'h3E71F996,
32'h3E7C7CD5,
32'hBD498566,
32'hBDC78B32,
32'hBD67FAB4,
32'h3ED536E5,
32'hBFCC0A36,
32'h3EA06D48,
32'h3DA0CAAD,
32'h3F0E3127,
32'hBEDAF7AB,
32'hBDC5B9F1,
32'hBD3C99C5,
32'h3D20B138,
32'hBE07BD76,
32'h3E3047D9,
32'h3E110397,
32'hBF989D91,
32'hBC8F2DD5,
32'h3F535A18,
32'hBE08241A,
32'h3EB483BB,
32'h3E162700,
32'h3E997E13,
32'h3CA64D6A,
32'h3E922A65,
32'hBC7C5D15,
32'hBD4DB46F,
32'h3E9AE6DE,
32'h3E264B0E,
32'h3E62080D,
32'h3EC8DD16,
32'h3E7EE9E2,
32'hBE6DF652,
32'hBD3E59B1,
32'h3E8E05B5,
32'hBF931A01,
32'hBC66C72F,
32'h3EC09130,
32'h3E5C94FD,
32'hBE91858F,
32'hBC91DDCE,
32'hBE4DA906,
32'hBD32232E,
32'hBE0B79CA,
32'h3EBE50A7,
32'h3ECE3149,
32'hBFA83574,
32'h3D41AA85,
32'h3F0ADA50,
32'hBDF2A474,
32'h3EA85AE7,
32'h3F0B5DF7,
32'h3E3B0836,
32'h3EAC89A0,
32'hBE117956,
32'hBD50FFE0,
32'h3D3630DC,
32'h3F28DF09,
32'h3DDF4C40,
32'h3CE18A33,
32'h3F2322D0,
32'h3EDA7481,
32'hBE5D4AFA,
32'hBE709701,
32'hBDBFCE75,
32'hBF37CC16,
32'h3E5389CD,
32'h3EEC2F86,
32'h3F169734,
32'hBF081AE3,
32'hBE472BCD,
32'hBD51615D,
32'hBC2627A1,
32'hBCEB602B,
32'h3EA8E5E5,
32'h3F05A356,
32'hBDCA9811,
32'h3E9EB801,
32'h3D3A938C,
32'h3E6B6B2E,
32'h3E947F23,
32'h3F282691,
32'h3E849A37,
32'h3D81B4F6,
32'hBE70A328,
32'hBCDB6C75,
32'h3CECCBA9,
32'h3EE3A02A,
32'h3DF9FA9E,
32'h3DFFF821,
32'h3F284D2C,
32'h3EF1DAF3,
32'hBE38FCCF,
32'h0EDD4862,
32'hBE64F076,
32'hBDB6FE63,
32'h3EA07F36,
32'h3F2FF8E7,
32'h3F355592,
32'hBE8D574F,
32'hBE4526FC,
32'hBCBD92E1,
32'hBC8FDABD,
32'hBE502214,
32'h3E5C6F55,
32'h3EAFDA6D,
32'h3E79A861,
32'h3EDBFBC4,
32'hBE6D5182,
32'h3EC98C93,
32'h2EC58AF0,
32'h3EDF7315,
32'h3EFCAAA8,
32'hBE8B08C2,
32'h3D7BC089,
32'h2EC9C2A8,
32'hBD5F1EBE,
32'h3EA428FC,
32'hBDC7EA6A,
32'h3E3387C7,
32'h3F05BBF9,
32'h3E9B58CB,
32'hBED4F2CF,
32'h3E1D997E,
32'hBEA8F5D0,
32'hBEECB149,
32'h3ECDDE09,
32'h3F40ABE8,
32'h3F28DC62,
32'hBEDBEC6C,
32'hBDDD6A58,
32'h3E538660,
32'h3EB20D1F,
32'hBEB3856D,
32'h3E53FE43,
32'h3E1EAF48,
32'h3E498F3E,
32'h3F031971,
32'hBE603E03,
32'hBD47CFC5,
32'h3E0A7AB1,
32'h3DF0FB8A,
32'h3E5A1722,
32'hBE517A64,
32'h3EB69478,
32'hBE11D028,
32'hBCD0C47A,
32'h3EA54703,
32'h5DEAE165,
32'h3EB66892,
32'h3EB4BC19,
32'h3DACC635,
32'hBDEA2C06,
32'hBE29D552,
32'h3D814C5C,
32'hBE9B7BDB,
32'h3E8491ED,
32'hBCDF6B07,
32'h3E8EFE13,
32'hBE212B2C,
32'hBDEE1669,
32'h3E042BC7,
32'h3EDA093B,
32'hBE9A0303,
32'h3E662CEC,
32'hBEF6B939,
32'h3EEC03C9,
32'h3E883476,
32'h2EC55EE8,
32'hBEE605B4,
32'h3EB07352,
32'h3DBC86F4,
32'hBD397CA8,
32'h3D792FAA,
32'h3EE8D934,
32'hBD487C0D,
32'h1DCDD5B9,
32'h3EF42618,
32'h3DA4DFC6,
32'h3E77221D,
32'h3D227E89,
32'hBEB92348,
32'hBD0ED0D5,
32'h3E87D354,
32'h3E4E6854,
32'hBD4225A4,
32'hBDB59D88,
32'h3CECC13A,
32'h3E6A1CD8,
32'h3E02B9C3,
32'h3E25489A,
32'hBEC4603F,
32'hBDBA3AF6,
32'hBF0BF3CA,
32'h3DEDD753,
32'hBEE68533,
32'hBDEE311C,
32'hBCCAFD1D,
32'hBE02E305,
32'hBE95B826,
32'h3E03A9C3,
32'hBE08CBDF,
32'h3D9249D4,
32'hBDEFFA18,
32'h3DD7B07B,
32'hBD9659DE,
32'hBC254325,
32'h3E1EB4C3,
32'h3EAB614A,
32'h3D4FF524,
32'hBD8AEF10,
32'hBF2E9065,
32'hBD7D2C37,
32'h3E5F382E,
32'h3E62D077,
32'hBE1E5530,
32'h3DC8EA24,
32'h3EB838DA,
32'h3C949E91,
32'hBD1F343C,
32'hBE16E2AB,
32'hBD25E350,
32'h3E9D5F27,
32'hBE74F90D,
32'h3E89522C,
32'hBF1F3248,
32'hBDB9D1FC,
32'hBDE62EF5,
32'hBD98753C,
32'hBE535D91,
32'h3E165CF7,
32'hBDF3A249,
32'h3CBB8BDD,
32'h3E0D05E7,
32'h175D1B98,
32'hBD26D2CF,
32'h3CD0C6A4,
32'h3E143FB0,
32'h3E476EBE,
32'hBE025466,
32'hBDF58193,
32'hBCF83D56,
32'hBCEC4D67,
32'hBDCCAD45,
32'h3E7FC1EF,
32'hBE95F933,
32'h3E29EBF7,
32'h3E3C28CA,
32'h3E0465B6,
32'h3D308B80,
32'hBEDCD574,
32'h3D9546EC,
32'h3ED19136,
32'hBDFF96FD,
32'h1DE6FB2F,
32'h3EB31C81,
32'h3D68FA80,
32'hBE13319D,
32'h3DADA0C5,
32'hBE415E77,
32'hBDF251AC,
32'h3E1D8CF2,
32'h3D8E1DAF,
32'h3E39B93A,
32'hBDA6CE63,
32'hBD430791,
32'h3D93B7D4,
32'h3E006DF2,
32'h2ED6F5E4,
32'hBD28DFF9,
32'hBE015B7D,
32'h3E7CFCD3,
32'hBE07BE08,
32'h3C1018DF,
32'hBD3C6C23,
32'hBEB7A238,
32'h3E238AB6,
32'h3DC3966E,
32'h3E989A85,
32'h3E066A53,
32'hBE6225CA,
32'h3E325199,
32'h3E600B05,
32'h3E259A95,
32'hBD409772,
32'hBF8125BB,
32'h3E2C7580,
32'h3DD03386,
32'hBDA0330C,
32'hBF430D84,
32'h3D96BF63,
32'h3E9E4725,
32'hBE4DCA00,
32'h3C54A14D,
32'h3E644E0F,
32'h3C89357E,
32'hBD7F9F13,
32'hBDEB27F1,
32'h3E65B76D,
32'h3E18D837,
32'hBE95D20A,
32'h3F1C4B8E,
32'hBDEB5235,
32'hBEE13022,
32'h3E4EF100,
32'hBF0C897D,
32'h3DA9B2CE,
32'h3EBC12F9,
32'h3E6F509E,
32'h3E02B7F3,
32'hBF2D8124,
32'h3E989CD9,
32'h3E929384,
32'h3DEACB81,
32'hBE4BC42A,
32'h3E88F55E,
32'h3D1FAFD3,
32'h3E78D580,
32'hBDF14245,
32'hBEC40314,
32'hBE3EFC73,
32'h3EC30FD1,
32'hBEC3F5A5,
32'h3DD39ABB,
32'h3E2B41AC,
32'h3D27F67E,
32'h3D168278,
32'h3DF26668,
32'h3D3F60B4,
32'h3D21C9F6,
32'hBE1A44C7,
32'h3DF5CA69,
32'h5DDF3538,
32'h3E42FAB1,
32'hBC8129F1,
32'hBF590CA7,
32'h3C54C27C,
32'hBE56397E,
32'h3E3AB4B3,
32'h3D5BE415,
32'h3E741D1B,
32'h3EB1CD5C,
32'h3D87E16F,
32'hBD1C8CE6,
32'h3D659334,
32'hBEE682BD,
32'h3DB0872C,
32'h3CC0FD8A,
32'h3D7E5E62,
32'hBDD4D52F,
32'h3E033FE7,
32'h3E38D382,
32'hBECA7F34,
32'hBD405125,
32'hBE8316CD,
32'hBDE7389C,
32'hBD1DDF6E,
32'h3E9422E0,
32'h3D8E5792,
32'hBE3A02B3,
32'hBE6C2C3C,
32'h3E923F1F,
32'hBD75E24F,
32'hBE8A9E56,
32'hBE8FD46B,
32'hBF4E201D,
32'h3C8106F1,
32'hBE283101,
32'h3E5E39D7,
32'h3DC420A2,
32'hBE6B73CB,
32'h3D69549E,
32'h3DD21EA8,
32'h2ECC1161,
32'hBE03C9A5,
32'h1DE8AFB3,
32'hBEEE12A1,
32'hBDFE6260,
32'h3E8D745E,
32'h3DDD058B,
32'h3DFF35DD,
32'h3EBA48E2,
32'hBF5E3467,
32'h3EF51EEB,
32'h3EC5183E,
32'h5DCA1DBF,
32'hBCEC6025,
32'h3D53B7A7,
32'h3E1B6186,
32'h3D1FA244,
32'hBE5AE227,
32'h3EFBD427,
32'hC0E00010,
32'hBEBB039C,
32'h3CD6F2CA,
32'hBF895AA5,
32'h3DD1DCA8,
32'hBE4E5F4B,
32'h3E57DCF6,
32'h3E9EE732,
32'hBF55D079,
32'h3DA11EB6,
32'hBEC92676,
32'h3D8BAF9E,
32'h3E1A6EA6,
32'hBEE6374B,
32'hBE882834,
32'hBE4AB367,
32'h3F140484,
32'h3E002486,
32'h3EB90975,
32'h3EAF4D84,
32'hBF4116F5,
32'h3F5DCE3E,
32'hBDB91588,
32'h3D24C424,
32'h5DD140D7,
32'h3D4F855D,
32'h3C9E24F2,
32'hBE8B17FE,
32'hBDBA72BB,
32'h3EAAD076,
32'h3E9E24EC,
32'hBF05F4BB,
32'hBF1FC156,
32'hC00F77BB,
32'hBC131E1C,
32'h3E886126,
32'h3E391367,
32'h3E6D728B,
32'hBF7F2D60,
32'h3E7E92DA,
32'hBE2C970A,
32'h3D503B20,
32'hBF17C292,
32'hBEE5EB24,
32'hBF8BD742,
32'hBEAA44DB,
32'hBE09955B,
32'hBEC573E8,
32'h3EB6AADC,
32'h3EC4EBCE,
32'h3D67E8BA,
32'h3F028A3A,
32'h3E28C4CD,
32'hBDFFD904,
32'hBD4E5138,
32'hBE811D17,
32'hBE824490,
32'hBDF356C8,
32'hBDBED1C7,
32'h3D5C665A,
32'h3E451EBF,
32'hBF14053C,
32'h3DC17FAB,
32'hBF9FFF21,
32'h3DAE4B86,
32'h3E8EA085,
32'hBE0EF677,
32'h3C2696CB,
32'hBD871A2D,
32'h3E531F8E,
32'h3EADE4E0,
32'h3E960677,
32'hBE7F738D,
32'hBC9FB801,
32'hBF949EE4,
32'hBF05AD69,
32'hBDF963B5,
32'hBF3461E6,
32'h3F9DB2F2,
32'h3CBC9D78,
32'h3ED7EB78,
32'h3E024149,
32'hBEDE3AA9,
32'h3D1BF955,
32'hBC77BDA4,
32'hBE8960F0,
32'hBEACB089,
32'h3E9DEB2A,
32'hBD95B358,
32'h3F35F85B,
32'h3EA7919D,
32'hBF4AB1D1,
32'hBE8B39B7,
32'hBF57B6D3,
32'h3DE3750E,
32'hBFBFC19C,
32'hBCB597BD,
32'hBF1B174C,
32'h3E23B946,
32'h3DE6F663,
32'hBF12012B,
32'h3EEA69CB,
32'hBDCB78F4,
32'h3F629054,
32'hBE4EDC14,
32'h3F52FF5A,
32'hBF3D9791,
32'hBC19A1DF,
32'h3F64A9BB,
32'h3C749D8A,
32'hBA4F7B9,
32'h3DE7A757,
32'hBEC1DDA3,
32'hBC439B06,
32'h3CE6D278,
32'h0EC49FA5,
32'hBE266A2F,
32'h3F549914,
32'h175BD240,
32'h3F053AB2,
32'hBF83ECA3,
32'h3E6E12F2,
32'hBF3FA65E,
32'hBF516BB4,
32'hBEC44EA8,
32'hBE2ABAC3,
32'h3DB37360,
32'hBE93D754,
32'h3E04F54F,
32'h3DE09763,
32'hBF2617E2,
32'h3E34365D,
32'hBE60ADBE,
32'h3F15F171,
32'h3D0BA7B1,
32'h3FC2C168,
32'hBF3313BC,
32'h0ED5EB9D,
32'h3C532D1B,
32'h3F1CA9DB,
32'h3E7849F6,
32'h3F5DC515,
32'h3E727E6C,
32'hBD1D65EB,
32'h3D9B4E3A,
32'hBECE86A5,
32'h3EE0D73B,
32'h3E8BA049,
32'h3D9C0475,
32'h3FC638DB,
32'h3D08292C,
32'h3D0A32FD,
32'hBE9435D4,
32'h3EFA7605,
32'hBF20B044,
32'hBEB0B27B,
32'hBF6E6F9E,
32'h3F70B74F,
32'h3E897C55,
32'h3F7BA777,
32'h3E7E04C3,
32'h3F95D0E7,
32'hBF2072BE,
32'h3C0FC770,
32'hBD40ED34,
32'hBDA967AD,
32'hBE682201,
32'hBCCA0CA3,
32'hBE24E1DA,
32'h3F3F6506,
32'h3D6DE811,
32'h3D80D47E,
32'h3E015E05,
32'h1DF762A4,
32'hBCCBE129,
32'hBE395C6C,
32'h3F41EF61,
32'h3C019F81,
32'hBE860070,
32'h3F4B95C4,
32'h3DAE8819,
32'h3C74F9AB,
32'h1DC134FF,
32'h3E12A1E0,
32'hBECF8D4A,
32'hBE52301F,
32'hBF3BB8EC,
32'h3EE96F44,
32'hBDB04E55,
32'h3F52CC92,
32'hBD63EA55,
32'h3D33033E,
32'hBED99CED,
32'hBD87E554,
32'hBD02AF8F,
32'hBDAEBFD5,
32'hBD344C7C,
32'hBDAB85F3,
32'hBD8B0697,
32'h3D85F9BC,
32'h5DE13AC8,
32'h3D5F8067,
32'h3CC87870,
32'hBC6C74EB,
32'h3D948532,
32'hBCF4C137,
32'hBD9EB3C1,
32'hBC822590,
32'hBD643753,
32'hBCAB4A4A,
32'h3D82634B,
32'h0EC5080E,
32'hBC8E85D8,
32'h3D9BF6BD,
32'h3D3BFE0C,
32'h3D07448A,
32'hBD90F4AA,
32'h3D4BD53E,
32'h3C801DEB,
32'h3D40E372,
32'h3DAAC2D4,
32'hBC33CEEA,
32'h1DEB58A5,
32'hBCAEAF8B,
32'hBC0685DC,
32'h3E56C109,
32'h3D7A96CF,
32'hBD366253,
32'hBE9DAAD9,
32'h3E5F9CB9,
32'hBDC32266,
32'h5DD00FB7,
32'h3DA35A5B,
32'hBCDCF4F3,
32'hBD1649C6,
32'hBEC19932,
32'h3E8B07F5,
32'h3E9123D1,
32'h3DABE559,
32'hBCB7F196,
32'h3D045A02,
32'h3E9CD33C,
32'h3CE427A7,
32'h3E183D3B,
32'h3EE8BA49,
32'h3D26DB48,
32'hBD89CC49,
32'h3DC49230,
32'h3D341AC0,
32'hBCDE5ACF,
32'h3D5783C2,
32'h3D32688A,
32'hBE16A6EE,
32'h3E181064,
32'h3F5AB59C,
32'h3E31D0FF,
32'h3F6301AA,
32'hBECCF29C,
32'h3FBF5CC4,
32'hBE51DC7B,
32'hBDA85D75,
32'hBE15B782,
32'hBEC7A426,
32'h3D490342,
32'h3CA392A6,
32'hBEDDF3F7,
32'h3EFA8268,
32'hBDCF1115,
32'h3E2B54AA,
32'hBDBDBEFA,
32'h3F125872,
32'h3E31ADE3,
32'h3E24048F,
32'hBF133809,
32'h3F0230B6,
32'h3CDF74C9,
32'hBE07FB06,
32'hBF1F9AB5,
32'h3F69AA2A,
32'hBD9EAD04,
32'h3C42CB41,
32'hBDAF08D4,
32'h3E3C563C,
32'hBE296027,
32'hBF5576DC,
32'h3DA1CE18,
32'hBD815C43,
32'hBEB3504A,
32'h3C653C8B,
32'h3D687DD5,
32'h3F291946,
32'h3EACB38E,
32'hBEC14044,
32'hBCAB6BAC,
32'h3CE97BF4,
32'h3DBE052B,
32'h3E106210,
32'h3D29A78D,
32'h3D0C7C1B,
32'h3DE8EA35,
32'h3D01EC66,
32'hBE06D295,
32'h3F0A73CA,
32'hBE5F31A0,
32'h3E305B99,
32'hBEBF534B,
32'hBE86788E,
32'h3F6F5245,
32'h3CCF7F9B,
32'h3EFA0C20,
32'hBE07DA34,
32'hBD19F956,
32'h3E6D59AD,
32'h3F180251,
32'hBF1CE9CB,
32'hBCF01949,
32'hBCDD445D,
32'hBF5B896F,
32'hBDD4F8AB,
32'h3D1CEE71,
32'h3D3A9094,
32'h3E40A23C,
32'hBF23D0E1,
32'hBD670B4B,
32'hBD0604E3,
32'h3F00EA48,
32'h075FF319,
32'hBD456B1C,
32'hBE116F08,
32'hBCD4ACED,
32'hBF6AF198,
32'hBFCCD2AA,
32'h3CEBC83E,
32'h3EA58FA2,
32'hBE24C28E,
32'hBF6DC9E9,
32'h2E4CD82,
32'h3E95749B,
32'hBEAF3991,
32'h5DC8D9AE,
32'h3EDCE705,
32'hBD504D81,
32'hBE4E5B8A,
32'hBEA97CA7,
32'hBEAA62C9,
32'h3EAD45DF,
32'h3DCC8DD9,
32'hBF0044BB,
32'h3E20E535,
32'h3E24BAA6,
32'hBE1EF22D,
32'h3DEF1625,
32'hBFAE874F,
32'h1CF618E,
32'hBD3E9EFD,
32'h3E307A77,
32'h3EB1E951,
32'h3E357611,
32'hBE497973,
32'h3EABA403,
32'hBEA9CDD1,
32'hBEF5458A,
32'hBD44553A,
32'h3DF65709,
32'hBE4ABC41,
32'hBF2BDE69,
32'h3D894271,
32'h3EEF0706,
32'hBF0A4BEB,
32'h3DA17361,
32'h3E6DFDC5,
32'h3EF22C0D,
32'hBF37F4D3,
32'hBC394051,
32'hBF2AE80B,
32'h3E3D6011,
32'h5DCB1F9A,
32'hBF1F00C8,
32'hBE3E1D19,
32'h3C580B10,
32'hBDDF046E,
32'hBD528C44,
32'hBF487014,
32'hBD11EAC6,
32'hBC805210,
32'hBE5802E8,
32'h3CF85387,
32'h3DDCD6A5,
32'hBC6032F8,
32'hBEAD7F9C,
32'hBEC6FDF8,
32'hBEAB5342,
32'h3E00A89D,
32'hBFFEF3D1,
32'h3E9F32E6,
32'h3E33C060,
32'hBD67E705,
32'h3DF3F492,
32'h3F18D326,
32'h3E7A5B73,
32'h3EE84984,
32'hBED06139,
32'h3C0C86ED,
32'h3E01772E,
32'hBF63D5B1,
32'h3DBB66CF,
32'h3DF0BEAC,
32'hBE3D0451,
32'hBE17BD46,
32'h3DBB4CA2,
32'hBDE3324D,
32'hBDDD59F6,
32'hBF211EB9,
32'h3C61791C,
32'hBDCA677A,
32'h1DE600F2,
32'h3E898090,
32'h3E25D305,
32'h3D0BD2A7,
32'h3E73FC18,
32'hBEABA944,
32'hBF25DD5E,
32'h3E3A6562,
32'hBFBCD198,
32'h3DBF60E6,
32'hBC763771,
32'h3C512F49,
32'hBDBBD25C,
32'h3F402AEE,
32'h3E9D4E74,
32'h3E617F57,
32'hBE2165CE,
32'hBD85B66A,
32'h3E081E9C,
32'hBF755486,
32'h3EA72088,
32'hBC420E2C,
32'h3E3F66DF,
32'h3DDDF812,
32'h3C5C1101,
32'h2E403C1,
32'hBE73A59C,
32'hBEF47B1A,
32'h3C6F71BF,
32'h3D1D5FC4,
32'h3C1845AF,
32'h3EBB8A48,
32'h3F054E2B,
32'hBD214004,
32'h3D78751E,
32'hBEF97895,
32'hBF8EE36E,
32'h2ECEB462,
32'hBE9FB5EC,
32'h3DD44B73,
32'h3D034586,
32'h3E397E23,
32'h3DEFC36D,
32'hBC0AD7E5,
32'h3E8E4F5A,
32'h3E383370,
32'hBE37ACDC,
32'hBE51ECF2,
32'h3E18DC7F,
32'hBFBA92F2,
32'hBDD41715,
32'h3F0387DA,
32'h3C4BAE5A,
32'h3E9D22B6,
32'h3D9C1C38,
32'h5DF02A18,
32'hBE6E3DE4,
32'h3EE65B8C,
32'hBE0CCFE8,
32'hBDECFBB7,
32'h3CEA9FDA,
32'h3E931F41,
32'h3DFBF2FE,
32'hBD9A0BC4,
32'h3DB8DD36,
32'hBF5039E9,
32'hBF447F28,
32'hBF19788F,
32'h3F1D4096,
32'h3CFE325A,
32'hBE2251EC,
32'h3E5EDA04,
32'h3DC7F088,
32'hBE883F1A,
32'h3E428F37,
32'hBD4EA7DD,
32'hBE1C1320,
32'h3D9CD555,
32'h3E1D5A05,
32'hBCB775FB,
32'h3DAB2BC5,
32'h3EE8C993,
32'h3D686C9D,
32'h3EC708B1,
32'h3D2399A2,
32'h3D3685B9,
32'h3E44B18E,
32'hBE65EDE0,
32'hBDD689A3,
32'hBD02721A,
32'h3EDEFD6B,
32'h3DF7B3C3,
32'h3DDAC088,
32'h3C4A1F48,
32'h3E23F2AE,
32'hBE69488A,
32'hBF812A0D,
32'hBED1875F,
32'h5DCB0B06,
32'h3DC13E9D,
32'hBC245669,
32'h3E8580D5,
32'hBDEEC2AB,
32'hBE7D1F39,
32'h3E4177F7,
32'h3E09E09E,
32'h3E1FAC33,
32'h3EB0B59D,
32'h3ED96371,
32'h3CB94830,
32'h3ED85A48,
32'h3ED5334C,
32'h3E8E84EB,
32'h3E5DF072,
32'hBD473BDB,
32'h3DD02C7D,
32'h3E1D788B,
32'h3C8B726B,
32'hBDCEDC58,
32'h3D392FE1,
32'h3EEA69E3,
32'h3E311CA2,
32'h3DD90FB7,
32'hBD12CD5F,
32'h3DA7810C,
32'hBE9691F8,
32'hBEE54AF2,
32'hBEAFFC27,
32'h075B5B64,
32'h3E9C883F,
32'h3EA424B7,
32'h3E95F6A7,
32'hBE96F8B5,
32'hBD15886C,
32'h3E7A474B,
32'h3E3E6D25,
32'h3DFD1A99,
32'h3DE6034C,
32'h3E963026,
32'hBE71B533,
32'h3EA5AD32,
32'h3E4C9CBB,
32'h3E12EA34,
32'h3CBE5CA8,
32'h3CEC1B86,
32'hBCE2ABF1,
32'h3DEC5D77,
32'h3EE3FC2C,
32'hBD586B56,
32'h3C5006E4,
32'h3EB1D2DB,
32'hBDDF5243,
32'h3E0585E5,
32'h3C201928,
32'h3D626E12,
32'hBD858093,
32'hBE6B1BF8,
32'hBE3FAB21,
32'h3DD4D461,
32'h3DC94BD6,
32'h3E5F2173,
32'h3EBF1818,
32'hBE269A94,
32'h3C907508,
32'h3D2D4434,
32'h3DE8F131,
32'hBEB95656,
32'h3EBDF086,
32'hBE90466E,
32'h3E867418,
32'h3E19FDEA,
32'h3D7ED3C2,
32'hBD90F55E,
32'hBD71BFA2,
32'h3E34C8DC,
32'h3EA80A76,
32'hBE91C2EA,
32'h3E28A5E2,
32'hBD9033BD,
32'hBD71C6BE,
32'h3E4922CF,
32'hBEC5E3E3,
32'h3D73BF5B,
32'h3DBF63D7,
32'h3D235FF5,
32'h3E3ADB75,
32'hBE5819C6,
32'hBE056E8B,
32'h3D4F4E06,
32'h3E985BC8,
32'h3F14C444,
32'h3E2C8903,
32'hBE506C67,
32'hBEA2D717,
32'hBD0C3142,
32'h1DE33821,
32'hBED8CE58,
32'h3EE55C43,
32'hBEDF2544,
32'h3ECA7AD2,
32'h3CEFFC38,
32'hBE30F161,
32'hBF038559,
32'h3DE6CD6D,
32'h3D4B7160,
32'h3D9A270D,
32'hBE8315A3,
32'h3E325EAE,
32'hBCCED8FE,
32'h3D7CB1A1,
32'h3E9FC2A5,
32'hBE0D6F0F,
32'h3E543DF5,
32'hBE41499A,
32'hBDA9131B,
32'hBDBFC510,
32'hBD499E4F,
32'h1DC63821,
32'h3E6DD78C,
32'h3D4CFBDF,
32'h3EA08901,
32'hBE1B77A3,
32'hBD7F1721,
32'h3E88E746,
32'h3CCFDF49,
32'hBE0E9E6D,
32'hBF5F6DC9,
32'h3EDCB7D5,
32'hBF14C7BC,
32'hBDA8E84D,
32'hBCA87A8E,
32'hBDF496FF,
32'hBF2097BA,
32'hBD5161C6,
32'hBDB88D32,
32'h3DC9206A,
32'hBED56EC1,
32'h3CEF0B03,
32'hBCFFFE5F,
32'hBD5C9B75,
32'hBD2FCB03,
32'hBD056BDE,
32'h3E2F55DF,
32'hBDAB02C6,
32'h3E93797E,
32'h3C644156,
32'hBEC97C4E,
32'h3E6149D5,
32'hBE7DF3BF,
32'h3E5A41D0,
32'h3EC90C42,
32'h3C9967AA,
32'hBDAEAAD4,
32'h3D484177,
32'h3EB4CBDB,
32'hBD53507C,
32'hBF3F055B,
32'h3E708D73,
32'hBF1A4ED7,
32'h3CC2249A,
32'h3D035729,
32'hBDAD1572,
32'hBF199BE7,
32'h3D9C90D7,
32'hBE103B38,
32'h3C10191D,
32'hBEB12F3F,
32'h3EA348BC,
32'hBC5C172F,
32'h2EDB08DC,
32'hBDD06149,
32'h3E71EEE8,
32'h3E83EBBB,
32'h3DAAF4EE,
32'h3E58B5A7,
32'h17596A57,
32'h3D23E9D1,
32'hBD1550F6,
32'hBD469021,
32'h3E2C268F,
32'h3C93B9FE,
32'hBD0945A2,
32'hBDB63EB8,
32'hBE9BAD76,
32'h3E444CEB,
32'h3E60B1A0,
32'hBEDC2162,
32'h3D88E59F,
32'hBDA93533,
32'hBD909CE3,
32'hBCED6D9C,
32'h3E444BE8,
32'hBF72A92E,
32'h3E9A84FE,
32'hBE652569,
32'hBE9DD1C1,
32'hBF0B4875,
32'h3E0B45BB,
32'hBD582B38,
32'hBDE16CF6,
32'hBC044E3B,
32'hBD8B80F9,
32'hBE024D75,
32'h3D834B7D,
32'h3E8C1833,
32'h3C354ABC,
32'hBEED227A,
32'h3DE29C72,
32'hBEB8DB94,
32'h3DCD97F0,
32'h3D803947,
32'hBE327354,
32'hBE6B3D8E,
32'hBE9192C9,
32'h3E42DBA8,
32'hBE60FE74,
32'hBE233EC7,
32'hBD74CAFC,
32'hBF2F34C2,
32'hBD344084,
32'hBD4DF1BE,
32'hBD7E5949,
32'hBF19A93B,
32'h3E46EDEF,
32'h3D8C7F15,
32'hBE72F86C,
32'hBEB8C2C6,
32'h3EADC5AB,
32'hBD04DFDF,
32'hBD78472E,
32'h3D0C5B9D,
32'h3DD39E56,
32'hBE6B7B42,
32'hBC5EF042,
32'h3D23DF4C,
32'h3D76D6E7,
32'hBED5B7F9,
32'h3EE97A75,
32'hBE5D9B39,
32'hBC3CA450,
32'h3E5268E3,
32'hBE6F7E84,
32'h3E830A78,
32'hBF9B6E49,
32'h3DCEB350,
32'hBD414BD8,
32'hBE986B64,
32'h3D94132D,
32'hBEB22D39,
32'hBE65CC87,
32'h3CC90649,
32'hBE776F49,
32'hBCB8495D,
32'hBE27CA8D,
32'hBE04668B,
32'hBECBDEB9,
32'hBEB2D78E,
32'h3DB07992,
32'h3CA648D8,
32'hBD2C29BC,
32'hBDB1AEC1,
32'h3DFBECD4,
32'hBCCEF55A,
32'hBDBF8498,
32'hBC39C961,
32'h3E3652F6,
32'hBEC57755,
32'h3E689388,
32'hBF0C3748,
32'hBE2E9E22,
32'h3E5C13C4,
32'hBE2B158E,
32'hBE0FA462,
32'hBF35C7C2,
32'h3E5C7D89,
32'h3E1F727B,
32'hBE59AB7B,
32'h3E2288B3,
32'hBFFCE1E1,
32'hBF07EFB7,
32'h3E34DDBA,
32'hBED37A52,
32'h3DE98A9E,
32'hBE539348,
32'hBD224661,
32'hBEEC21EF,
32'h3E3B6A3A,
32'hBE095D93,
32'h3C42ACF3,
32'hBDB8D7B7,
32'hBDB76DA1,
32'h3D1B11F9,
32'h3EB6C695,
32'h0ED95B33,
32'hBDFB61ED,
32'h3E26336D,
32'hBF469EA0,
32'h3CEB3D5D,
32'hBF935F70,
32'h3E20BB66,
32'hBC9FD83A,
32'h07529390,
32'h3D624B5C,
32'hBFBFB866,
32'h3EEDB7C5,
32'h3CE9762E,
32'hBE3430F6,
32'h3DA7E580,
32'hBF3A5FC8,
32'hBF536B6C,
32'hBD43B4EC,
32'h1DDCF56E,
32'h3E193710,
32'h3EA9B1D0,
32'h3E722C98,
32'hBF4F306C,
32'h3E2F98E0,
32'hBCA84E1B,
32'h3D3A4906,
32'hBD10D230,
32'hBDCD8A1D,
32'hBEDA3493,
32'h3DEBC6FD,
32'h3E061DFA,
32'hBD7D94B1,
32'hBE0B004C,
32'hBF23712A,
32'h3E30D41B,
32'hBF6FAD43,
32'h3E6FF12F,
32'hBE51EFF5,
32'h3E5C3331,
32'hBD56679B,
32'hBF974823,
32'h3ED55AEB,
32'h3CC041D4,
32'hBE93E085,
32'hBE0DCBB6,
32'hBF05829A,
32'hBE14BE1E,
32'h3E09660B,
32'hBDD9C29B,
32'h3E4D1C5D,
32'hBD7D51BC,
32'h3ECF0E3A,
32'hBF054815,
32'h3E8E8C12,
32'hBE992071,
32'hBC290F8D,
32'hBD07E6BF,
32'hBE8A7C56,
32'hBEB37E20,
32'hBDA88568,
32'h3E4E0B0E,
32'h3EAF3657,
32'h3D8B19B6,
32'hBEBC58F4,
32'h3DEE7058,
32'hBF93FC90,
32'hBC8B6588,
32'h3D8B5EBC,
32'h3E7EDCD2,
32'hBF181B6A,
32'hBECF9F5B,
32'h3E9C2209,
32'h3D8DED52,
32'h3DCCF2DA,
32'hBF365F02,
32'h3E71C2E1,
32'hBEE573AC,
32'hBC968974,
32'hBDE12DAA,
32'h3DDF5546,
32'h3D9376D6,
32'hBEB03B93,
32'hBDCB13B3,
32'h3ECC4311,
32'h3E20DF7E,
32'hBDD733AC,
32'h2EC98151,
32'hBEFC8594,
32'h3D1B7C75,
32'h3ED0E662,
32'h3E3B34CF,
32'h3E382202,
32'h3DEA9E5E,
32'hBF7E07DC,
32'h3F2FA925,
32'hBE1B9C9C,
32'h3E858479,
32'h3F804490,
32'hBE7F6012,
32'hBF1427A7,
32'hBF0CD238,
32'h3E876E77,
32'h3F4174B0,
32'hBE662B65,
32'hBF4983F8,
32'h3F1635F1,
32'hBEAB0AA3,
32'hBEBAB638,
32'hBD5CD8D5,
32'hBEA5BD54,
32'h3FC211D5,
32'h3D35F6D1,
32'h5DD66E31,
32'h3E8A11FA,
32'h3DE272FE,
32'h3CEC1539,
32'h0ED38222,
32'hBE9843FA,
32'h3F166080,
32'h3F2BC4DE,
32'hBF0C19A0,
32'h3EDC00D1,
32'hBE3E5B46,
32'hBDA239A4,
32'h3F013A72,
32'hBEE1BA1B,
32'hBE3C83C1,
32'hBFA75501,
32'hBF042BFC,
32'hBEBB6314,
32'h17536B7D,
32'hBDAD8FAA,
32'hBEB9049B,
32'h3F49D39B,
32'hBF0F84C0,
32'h3F84FF6D,
32'hBE0CA2BA,
32'h3F9B868E,
32'hBE580374,
32'hBE9ACC32,
32'hBF0C4102,
32'h3F1E6B08,
32'hBD2BF2B4,
32'hBE4233AE,
32'hBEAB9623,
32'h17552F81,
32'hBCA0119B,
32'hBE821BFB,
32'h3E85CFF1,
32'h3F3C1A38,
32'hBE3E684C,
32'h3EFAD5F9,
32'hBEAFC164,
32'h3F4005F5,
32'h3C641655,
32'hBE6E3349,
32'h3E316995,
32'hBF83DC03,
32'h3EA1A76C,
32'hBEE9D4EA,
32'hBD9D4752,
32'h3EFA3BD7,
32'hBECEC9F8,
32'h3F0BD5CB,
32'hBE0B3D83,
32'h3F23EB19,
32'h3CD212EF,
32'h3FE93E4E,
32'h3F17B657,
32'hBDF1E91F,
32'h3E1E137F,
32'h3F1963D5,
32'hBD5DECF0,
32'h3FFC2A98,
32'hBC6EB2E1,
32'hBDBF4A25,
32'h3D73DF89,
32'h3F02A5F9,
32'h3FB79D17,
32'h3EBB6625,
32'hBEAF0720,
32'h3F908E0E,
32'h3DA6F729,
32'hBF3549BC,
32'hBF303589,
32'hBE6A49F1,
32'hBEAE71EC,
32'hBF2B8490,
32'hBF60997D,
32'h3FA047FA,
32'h3E81F01D,
32'h3EC41AD7,
32'hBD3E1503,
32'h3F3F10D6,
32'hBF15A68D,
32'h3C4E583E,
32'hBCF78F28,
32'h3CC1AFEA,
32'h3CC279F9,
32'h1DC1D449,
32'h2ECD658B,
32'h3C8A3574,
32'h3C80EB27,
32'h3D4748CD,
32'h1DF9AC7A,
32'hBD1FF37A,
32'h3DE81232,
32'hBD0EF8B2,
32'h3D44197F,
32'h3C9F9927,
32'h1DEA6602,
32'h5DE380C3,
32'hBA30F81,
32'hBD2F0ECF,
32'h3CFBF156,
32'hBE0F1C8C,
32'h3E653379,
32'hBD76937E,
32'hBD2B26F7,
32'hBC8B60AA,
32'h3CF9B14C,
32'h3EA8C7F6,
32'h3E09F259,
32'hBC0A7AB0,
32'h3DC9C0CD,
32'hBD566B38,
32'h3D64A6EB,
32'hBD84F513,
32'hBD8D6926,
32'hBD94F99C,
32'hBD58F63C,
32'h3C46D609,
32'h3DBF9260,
32'h3CAAF0E5,
32'h3D818F16,
32'hBD9A2ADE,
32'hBD5A3C60,
32'h3D8898AD,
32'h3CBDD0A2,
32'h3D1148C3,
32'h3DF2B5C2,
32'h2ED14937,
32'hBD0A3050,
32'hBD012FC5,
32'hBCE30373,
32'hBD477D8D,
32'h3D81A230,
32'hBD174790,
32'h2ED89E0E,
32'h1757FA1B,
32'h3C4B6C2D,
32'h3E0F6441,
32'hBD8EF445,
32'h3D61DAFE,
32'h3D2D4754,
32'hBDD5B664,
32'h3D89E7D0,
32'h3E22C1A6,
32'hBDCFDBA9,
32'h3CBC8ED8,
32'hBE82DC33,
32'h3E926751,
32'h3E41F0D8,
32'h3D3783C7,
32'h3D4C5766,
32'h3C1A3244,
32'h1757CB80,
32'hBEB8BCF7,
32'h3E8A198C,
32'h3EB6FD07,
32'h3ECD2B6E,
32'hBCCAEA1B,
32'h3D0F5978,
32'h3D68D97E,
32'h1DC4404B,
32'h3E146FFA,
32'h3F0DB231,
32'h3D43D804,
32'hBE233E58,
32'h3EC920E2,
32'hBC2A105F,
32'h3E30C942,
32'h3CF95158,
32'hBD8665EB,
32'h3D4DA653,
32'hBE214378,
32'h3E326BC0,
32'h3E5C740B,
32'hBE959B4D,
32'hBD3D7B4E,
32'hBF17730D,
32'h3E1925B0,
32'h3E364588,
32'h3F011A84,
32'hBDC8E08E,
32'hBCC8B366,
32'hBD131355,
32'hBF4487D5,
32'h3F5F38B6,
32'h3D971BE3,
32'h3DBE0559,
32'h3EDEDD4F,
32'h3EF68F0F,
32'h3D64072E,
32'h3DF012D2,
32'h3DAEFCE5,
32'h3F42516B,
32'h3DC3149F,
32'h3D25002F,
32'hBDD3F582,
32'h3C39442E,
32'hBF220F9E,
32'h3E74C643,
32'hBDC38E53,
32'hBDCF4625,
32'hBD707E97,
32'hBF94AE97,
32'hBF812D48,
32'hBF223316,
32'h3F03C2BE,
32'hBE931280,
32'hBD54BD09,
32'h3D79FFAB,
32'h3F293FFE,
32'h3D4C9F80,
32'hBCA1529D,
32'h3C0DB46C,
32'h3E4203BF,
32'h3F341078,
32'h3DB374E8,
32'hBEE9E83B,
32'h3F8116EA,
32'h3D8C6553,
32'hBF562515,
32'hBFA8C901,
32'hBE6A3CDD,
32'h3DD1CA3E,
32'hBE286F3B,
32'hBE95FD44,
32'h3F064E01,
32'hBF116F31,
32'h3DEAF946,
32'hBE91C823,
32'hBE6B5118,
32'hBE908034,
32'h3F11BDA4,
32'hBEF65280,
32'hBF185894,
32'h3EB158AD,
32'h3D8A9448,
32'h3EC2599B,
32'hBD8383D4,
32'hBE2A6D1E,
32'h3E73A922,
32'hBF88DA00,
32'h3D48C0E1,
32'hBD509E8F,
32'hBDEED721,
32'hBF10BDB0,
32'hBDA89C32,
32'h3DA66652,
32'hBE9D8EA0,
32'hBE5B3692,
32'hBFA9C04A,
32'h3E5DC970,
32'h3ED4BD7C,
32'h3E0B847A,
32'hBEE01DAF,
32'h3E8FB500,
32'h3DAD4531,
32'hBE5D7B52,
32'h3E2D64CF,
32'h3CA126B4,
32'hBEBF10A8,
32'hBF5BB3ED,
32'hBE271E2A,
32'hBE19ADBB,
32'hBD92F1C4,
32'h3D116E21,
32'h3DC42FE1,
32'h3ED3D696,
32'hBE11BEFF,
32'hBEBDEAC3,
32'h3D5C670E,
32'hBF37C155,
32'hBDCCD58D,
32'hBCF2742A,
32'h3EE60FA1,
32'hBD8AD7EE,
32'h3D96A821,
32'h3D07BFBE,
32'h3D9E48DB,
32'h3E60F77A,
32'hBF79B968,
32'hBF401A30,
32'hBF9933FE,
32'h3D06AB48,
32'hBED116FC,
32'h3CB44E50,
32'h3E7975D9,
32'hBF076599,
32'hBE6D58CF,
32'h3E8E7A7F,
32'h3C5DB5F2,
32'hBF3C1A8D,
32'hBE69D832,
32'hBF75B15F,
32'hBEC17646,
32'hBCCB8E57,
32'hBE449434,
32'h3EAB8CB2,
32'h3E76D579,
32'h3DCCFD56,
32'hBE022350,
32'hBF32BA39,
32'hBDF9C685,
32'hBD22DA36,
32'h3D4890FB,
32'hBE8128EF,
32'h3D2EAC4D,
32'h3E3C5960,
32'h0ED7BF78,
32'hBD708D6E,
32'hBF211CA4,
32'hBF68C0D6,
32'hC016ED74,
32'h3E81409A,
32'hBEAF10E5,
32'hBE3167AD,
32'h3F0FBC6E,
32'h5DEB3EDF,
32'h3E1A896C,
32'h3ED4F877,
32'h3D0F9C66,
32'hBF100A84,
32'h1750A882,
32'hBFD464C4,
32'hBD97AA08,
32'h3C89F733,
32'hBE95CA9E,
32'hBDAA9E48,
32'h3DAC95E8,
32'h1DF3460D,
32'hBE67227E,
32'h3F079CE5,
32'h3CC05CBA,
32'hBD9BB550,
32'hBE6471C2,
32'hBE698FBF,
32'hBDE4242D,
32'hBD4F3211,
32'h3EE2584A,
32'hBEB88822,
32'hBF2C9F3F,
32'hBE6B3CCC,
32'hBE3A02F3,
32'h3DECBB08,
32'hBE43731D,
32'hBE21571A,
32'h3DCCE476,
32'hBF23A4BE,
32'h3E36938A,
32'h3D923B7A,
32'hBE638094,
32'hBEB77AAB,
32'hBE28457B,
32'hBF7B914A,
32'hBDBE7BA8,
32'hBD3121EC,
32'h3E4E594C,
32'hBD252DBB,
32'hBD06B93E,
32'hBE069650,
32'hBCD43AAE,
32'hBE5C884D,
32'hBDA7B7DC,
32'hBD4E3BF4,
32'hBEEEC8CD,
32'hBDDEF605,
32'h3E16978F,
32'hBD8823B3,
32'hBE9D82D9,
32'hBE7F7736,
32'hBF80A715,
32'hBE951FAA,
32'h3F55CF6B,
32'h3E37E057,
32'hBDD701BA,
32'hBDB9B057,
32'hBD4141B8,
32'hBF2FF4FE,
32'h3DF1415C,
32'h3D4EAB36,
32'hBE498736,
32'h3DE2D767,
32'hBDCE7728,
32'h3E1089E5,
32'hBD374DFB,
32'h3DC3812E,
32'h3F006BB3,
32'h3DE3C1D6,
32'hBD92FBC5,
32'hBD7925C3,
32'h3DCC0F03,
32'h3E8519A3,
32'hBD67C58C,
32'hBD322E9F,
32'hBE509307,
32'h3D907DDE,
32'h3E70661E,
32'hBE1ABAFE,
32'h3E1B9100,
32'hBE77A8DB,
32'hBF68FBF9,
32'hBFA12053,
32'h3F141A12,
32'h3E1863E9,
32'hBD80AC13,
32'hBDE6C22C,
32'hBD58E383,
32'hBE8DE14C,
32'h3DFBC070,
32'h0755B329,
32'h5DE1578E,
32'hBE08B97A,
32'h3D968805,
32'hBDF3F40B,
32'h3E004096,
32'h3E8B83E3,
32'h3E588B73,
32'h3D7DA0D9,
32'hBD357BBD,
32'hBD9BBF6C,
32'h3DD3F2FA,
32'h3E4CBF06,
32'hBD6ACEC3,
32'h2ECEBF07,
32'h3DDFCFAF,
32'hBC9ED00C,
32'h3E4C3724,
32'hBD707871,
32'h5DCA9CCA,
32'hBE69CCA4,
32'hBF23D380,
32'hBF8F9E23,
32'h3E8AF7E9,
32'h2EDBEB84,
32'hBDD1E024,
32'hBECC4097,
32'h3E810634,
32'h3E1CFD68,
32'h3E0A8E49,
32'hBC766C8E,
32'h3E3B1932,
32'h3DA3C17C,
32'hBE555124,
32'h3D59A9CC,
32'h3CF9F288,
32'h3ECBE931,
32'h3C53A528,
32'h3D8CC19B,
32'h3DBB5733,
32'hBE2F6A0D,
32'hBE39039A,
32'h3C993CF5,
32'hBDD773F5,
32'h1DCBC9E9,
32'hBCBA677B,
32'hBD0B5323,
32'hBEE0EB62,
32'hBE29198C,
32'hBE400197,
32'hBE017D4E,
32'hBEF8EE81,
32'hBF1A790A,
32'h3E94B44A,
32'h07557415,
32'h075EE250,
32'hBCA23A8B,
32'hBE7932CA,
32'hBD9B8C51,
32'hBDC30848,
32'h3E0FF45D,
32'hBE1746AB,
32'h3E6E2E59,
32'hBCA40F3F,
32'hBD8D1A27,
32'h3DC2994E,
32'h3D4E45EE,
32'hBE858DA2,
32'hBE00ED1D,
32'h3E213BA3,
32'hBC0B1571,
32'h3D74936D,
32'h3E32A84A,
32'hBC1A99C9,
32'hBD823BA5,
32'h3DB6E4F1,
32'hBDA1F3A7,
32'hBEA42BAD,
32'hBE7CFA54,
32'hBD108315,
32'h3DCAFF2B,
32'hBE677915,
32'hBE1AB2A1,
32'hBDB2B08E,
32'hBDCD265B,
32'h3E51EF75,
32'hBEA33E7C,
32'h5DD82B58,
32'hBEBA0840,
32'hBE1199FF,
32'h3D1450EF,
32'hBE8BF052,
32'h3E9B6B0C,
32'hBE260622,
32'h3E0A7133,
32'h1DC42C08,
32'hBE29FFB2,
32'hBEA4A547,
32'h3D698A82,
32'h3E1F65E6,
32'hBD8135D4,
32'hBDEFAC99,
32'h3E4D7D3D,
32'hBC8D9863,
32'hBC6AFE84,
32'hBD8F6B44,
32'hBEC86D67,
32'h3DC4B55E,
32'hBE01D4C7,
32'hBE02D0F1,
32'h3D2965A8,
32'hBEA2B3F0,
32'hBD9C6509,
32'hBE407DF4,
32'h3ED6E94D,
32'h3F03F6A7,
32'hBCCEBC25,
32'h3DF43BA2,
32'hBE16AA3B,
32'h3D9E48B4,
32'h3D9D6F03,
32'hBEF003D0,
32'h3E8BB2AA,
32'hBEA4A45B,
32'hBD21064E,
32'h3DC95409,
32'h5DE32CFA,
32'hBFAFB366,
32'hBCA5A175,
32'h3E3DF9E0,
32'h3D5F7CE2,
32'hBE900B83,
32'hBDC29783,
32'hBDC78F15,
32'h3D33F735,
32'h2ED07B1C,
32'hBEB7C8D2,
32'h3DAF11C6,
32'hBDD6568F,
32'hBD9A2427,
32'h3D11BCFB,
32'hBEB2D148,
32'hBDD64E71,
32'hBE382334,
32'h3DC37A5C,
32'h3E937EE3,
32'h3C24EAC4,
32'h2E4E1A3,
32'hBCCE9031,
32'h3D8BFFF9,
32'hBE2543D7,
32'hBF6974B9,
32'h3C3B4A5C,
32'hBEF7118A,
32'hBEA7B8CD,
32'hBD8EF883,
32'h3DF32876,
32'hBF813446,
32'h3C2DAAD3,
32'hBCF004D9,
32'hBD4CFB2C,
32'hBE928BFB,
32'h3E5FB8F6,
32'hBD6F2D0F,
32'hBD3E4CDF,
32'hBD6D1E6A,
32'h3C95321A,
32'h3F03DB5D,
32'hBD8F0441,
32'h3DCD83E5,
32'h3E8E11AB,
32'hBEE8A7FC,
32'hBC593640,
32'hBE596486,
32'h1DFB33D5,
32'h3CE86765,
32'hBE066C0C,
32'hBD412889,
32'hBE676BC5,
32'h3E1F76FC,
32'hBC98B8F0,
32'hBF3BA075,
32'h3E53B36E,
32'hBF26DDA7,
32'h1CC1941,
32'hBCA1D994,
32'hBE60C1F4,
32'hBFDED06C,
32'h3E40774F,
32'h3DFBBF43,
32'hBE26C02F,
32'hBEBC36C8,
32'h3EA3D96D,
32'h075C309F,
32'h3DBB4663,
32'hBD0D6879,
32'h3CCCDB0A,
32'h3E8D1927,
32'hBDCC9FED,
32'h3D1C13B0,
32'hBE6D6511,
32'hBE6712A2,
32'hBDF14D55,
32'hBD1B73D9,
32'hBC0B1590,
32'h3E2ADAD0,
32'hBC60577C,
32'hBE888E35,
32'hBD9464B4,
32'h3E3B7004,
32'h3E1CB9B9,
32'hBF6A51C5,
32'h3E2DE42A,
32'h3DD33DD9,
32'h3E43B461,
32'h3E60357C,
32'hBE22D41E,
32'hBFD2FD60,
32'h3E784CB2,
32'hBE9C5B24,
32'hBDD55A27,
32'hBF1A125B,
32'hBEFBE0E1,
32'hBC88AFFB,
32'hBC95E7CB,
32'h3D6D2FD4,
32'hBE02ECE4,
32'h3EB10A36,
32'h3E4849C4,
32'h3DADB073,
32'h3E4B32A2,
32'hBEC0B627,
32'h3E7A106C,
32'hBE7F189E,
32'hBD4B8C49,
32'hBC999E0A,
32'h5DC5007A,
32'hBE8FB9C6,
32'hBE80BDC0,
32'h3E132660,
32'hBDEFE790,
32'hBF48C898,
32'h3E33B55A,
32'hBF3323C6,
32'h3D9F0196,
32'h3D540333,
32'hBEA1759D,
32'hBDE70482,
32'h3D9D787A,
32'hBD08086A,
32'hBDEEA8D4,
32'h3E1BC179,
32'h3E81A13A,
32'hBD70A914,
32'h3D19F069,
32'hBDD8C30C,
32'h3D60DE87,
32'hBD7BECF8,
32'h3E1E96C8,
32'h3D99643C,
32'hBC7496CA,
32'hBE93B63B,
32'h3E160655,
32'h3E103487,
32'h3DC55926,
32'hBC64897B,
32'hBDCD78BB,
32'hBDCB2F1C,
32'hBF3BAD49,
32'h3E45AFB4,
32'hBE1869F1,
32'hBE38E4B7,
32'h5DE26F17,
32'h3D904084,
32'h3D21C56F,
32'h3D619A59,
32'hBEDDFDA8,
32'hBE558455,
32'hBDF18921,
32'hBDA31DB4,
32'hBDDC26A9,
32'hBEE1A7AD,
32'h3D06B10D,
32'hBDFC8A48,
32'hBD3A0544,
32'hBF020BA5,
32'h3EBB5C80,
32'h3D8A22C0,
32'h3CF6B2EB,
32'h3EF7DE91,
32'hBDD4F379,
32'hBF1B2BFC,
32'hBE037F9B,
32'hBD0350AC,
32'hBDB9B407,
32'h3E1347D8,
32'hBD8C0766,
32'hBE3C3D02,
32'hBF7E7CB5,
32'h3E3C584D,
32'h3DD431AD,
32'h3E48A77D,
32'h3E967219,
32'hBF5D997C,
32'hBE772423,
32'h5DC8E92C,
32'hBEA7BDDC,
32'h3ED9D059,
32'hBDD82D13,
32'hBE32EC69,
32'hBE7F6CB5,
32'hBE62F62E,
32'h3E7C5DCC,
32'h3DFDDA92,
32'hBD97C4CE,
32'hBF182B9C,
32'h3EC70CAC,
32'h3E1F43C3,
32'hBD430847,
32'h3E5030F5,
32'h3F0EF33C,
32'hBF0F50E7,
32'h3EDCE3F9,
32'hBE3D23A1,
32'h3DF5BE19,
32'h3E9BA8FB,
32'hBC30EEC5,
32'h3DE2BFDB,
32'hBF771254,
32'h3DF83C82,
32'h3DF48638,
32'hBD01E62F,
32'hBF1AB396,
32'hBD4EA5F3,
32'hBCD74F30,
32'hBDE9E154,
32'hBEE68A17,
32'h3E96FBE1,
32'h3E2649D4,
32'hBED89E9C,
32'h3D859DAB,
32'hBE97521B,
32'h3E6A78C2,
32'h1DE21293,
32'h3D39948A,
32'hBEDA1B71,
32'h3F2BE778,
32'h3D814B5C,
32'hBDB8F4AA,
32'hBD35BA88,
32'hBE4DA603,
32'hBEF9F8D7,
32'h3EA3AC52,
32'hBF061FD5,
32'h3E180117,
32'hBE007845,
32'h3E3B6EC0,
32'h3CEA1643,
32'hBD350533,
32'hBDA64132,
32'hBE2BCACC,
32'h3E60B5BF,
32'hBF82273D,
32'h3EDEF930,
32'h3E16DE16,
32'h3EC5FF67,
32'hBE6EB26C,
32'hBDE595DA,
32'hBF44AFBD,
32'hBE9DC302,
32'hBE99B315,
32'hBF342CE2,
32'hBE18CA47,
32'hBD8D5A11,
32'hBD0A997B,
32'h3E160B29,
32'h3F181A96,
32'hBE000420,
32'hBE292A88,
32'h3F7E54AD,
32'h3E9C0D14,
32'hBF11589F,
32'h5DD336E1,
32'h3CF7C04B,
32'h3D1C0D65,
32'hBE13D9D2,
32'h3E2CAA55,
32'hBDCE6961,
32'hBE88E431,
32'h3E68F860,
32'hBD0C85DC,
32'h3EB34127,
32'hBF62DDAD,
32'h3ED8544E,
32'hBEB9E4F2,
32'h3F4D9DFF,
32'hBD10F904,
32'hBD8D7352,
32'hBF8C0654,
32'hBE30FB5F,
32'hBEBB3B48,
32'hBF1BC46B,
32'h3D1FC8E5,
32'h075CB461,
32'h3DEFB9D4,
32'hBEFACA70,
32'h3EC2134E,
32'hBE63853C,
32'hBECFB486,
32'h3DEDE45F,
32'hBE1362AE,
32'hBF83FB41,
32'h3EDFD493,
32'h3C1087EE,
32'h3EBC3FBF,
32'h3EEB8EA1,
32'hBEC20F7F,
32'hBE80A089,
32'hBF352F60,
32'h3F21507B,
32'h3F0B41F2,
32'hBDBDCCC5,
32'hBE90FBFD,
32'h3EE678CF,
32'h3F28D358,
32'h3EBD4B83,
32'hBDAF9317,
32'h3EC003B9,
32'hBE239EA0,
32'hBF10A6E1,
32'hBEF9B107,
32'hBEBF808F,
32'h3E2F8414,
32'h3C4C366D,
32'h3D763265,
32'hBF429785,
32'h3F1AFD4F,
32'h3F1C479E,
32'hBE8077DB,
32'h3F1ECFCD,
32'h3E99F171,
32'h3F059BE1,
32'h3F49844B,
32'hBEFDC9AC,
32'h5DC7F4F2,
32'hBFAAD0A7,
32'hBEE961A0,
32'h3EF691A6,
32'hBD8A774F,
32'h3E97754C,
32'hBE3F6B10,
32'h3E9729FE,
32'hBF65C807,
32'h3F35659F,
32'hBE203007,
32'h402FB346,
32'hBE49D9D3,
32'hBDBABCA6,
32'hBE2704F4,
32'h3F156F14,
32'hBE8D880D,
32'h3E839F9C,
32'h3F7E99A2,
32'hBD003DED,
32'h3D76B496,
32'h3D273510,
32'h3F147030,
32'h3F695FE3,
32'hBF8AFFA5,
32'h3FDB33A5,
32'hBE8DB88E,
32'h3F4C4867,
32'h3E4B0DB7,
32'hBE8BE12C,
32'h3D622A16,
32'hBEC342E2,
32'h3E3BEE48,
32'h3F69E725,
32'h3D3884BB,
32'h3ED9C08E,
32'hBF381F8F,
32'h3ED588E0,
32'hBF2A7D0B,
32'h3F662493,
32'h3D831BED,
32'h3F9387E2,
32'h3FCD7A67,
32'h0EDA42F0,
32'h3EEE0D1D,
32'hBC873233,
32'hBEE8AF26,
32'h3EAB2247,
32'h3F346BDF,
32'h3D2A73B6,
32'h5CEF330,
32'h3F436CAB,
32'hBEEFF227,
32'h3E2A0199,
32'hBF3B0E8F,
32'h3F929B02,
32'h3D20F4FB,
32'hBF920752,
32'hBED5E3B5,
32'h1DC61317,
32'h3F386981,
32'hBDBE2270,
32'h3EFCCAF2,
32'h3EC059F2,
32'h3D889DF2,
32'h3E13A3AF,
32'hBEBA62D3,
32'hBE055134,
32'h3EE62F96,
32'h3DE60B6B,
32'hBDBC712D,
32'hBD49B8ED,
32'hBD660BA8,
32'h3DB30BA5,
32'hBD4455BE,
32'hBD96F3BB,
32'hBD5B2D93,
32'h3D0DAB56,
32'h3D2F6040,
32'h3CE68D3D,
32'hBD4F1340,
32'h3CDBEEFB,
32'h3C1CFF65,
32'hBD3E4DF1,
32'h3D095C04,
32'h1DD6D141,
32'h5DDC96EF,
32'h3CB21432,
32'h3D0C4720,
32'hBDA36779,
32'h3C6C6DCC,
32'hBC9411F3,
32'h3C085C41,
32'hBCE5E981,
32'h3D641A65,
32'hBD9C97BA,
32'h3D910AD3,
32'h3D1B302A,
32'h075B274B,
32'hBCF5CCDF,
32'h3D90C006,
32'h3D327D83,
32'hBD9EDD9C,
32'h3D9E5639,
32'hBD6334B9,
32'h3D94F37B,
32'h3D0A2284,
32'h3D8171BE,
32'h3DD3A9C8,
32'h3DBEAA95,
32'h3C8561E5,
32'h3DCCEC6C,
32'h5DDD15FE,
32'h1DF1CFDB,
32'h3DD14D4B,
32'hBD918B6E,
32'h0ED7E759,
32'h3C46CEFD,
32'hBC93CFEB,
32'h3DB9E8A1,
32'h3DB23455,
32'hBDAB82C9,
32'hBCA3EB9F,
32'hBCC6C946,
32'hBC15A75B,
32'h3C1FDD7B,
32'h3C8DBB6F,
32'hBD88854F,
32'h3D32F6A2,
32'hBD8123C2,
32'h3DC991C1,
32'h3DA13B1F,
32'hBD345381,
32'h1DCC1934,
32'hBDEDB025,
32'h3E83B62A,
32'h3C56C5AB,
32'h3CC2E1B3,
32'h3CCE6E07,
32'hBD9E3938,
32'hBD9D359F,
32'hBC01AD8C,
32'hBDDF1425,
32'h3DC60A8C,
32'h3E5A55C3,
32'h3D52B853,
32'h3D8750BC,
32'h3CCF78A9,
32'hBC00C536,
32'h3D4FB771,
32'h3EDC90FD,
32'h3CB1969B,
32'hBD9FDE4B,
32'h3E82E086,
32'h3D5DCCB7,
32'h3E122F0B,
32'hBD8DC055,
32'h3C615FA5,
32'h3D710066,
32'h3E0097A7,
32'h3E40238F,
32'h3FC0ECB8,
32'h3D5C916D,
32'hBDFA8E66,
32'hBD978816,
32'hBD87BE2C,
32'hBE6CB3C3,
32'h3EB4A04C,
32'h075FF61D,
32'h1DC13D84,
32'h3CD5E6DC,
32'hBEC12346,
32'h3F2C33DA,
32'h3ED9C0CF,
32'hBE1056CD,
32'hBE3B7A47,
32'h3E0DA9E7,
32'hBE4B9704,
32'hBE8C5E16,
32'hBDBC5705,
32'h3EE70E83,
32'hBC7CB11F,
32'hBD6B65B4,
32'h2ED87DB3,
32'hBD332BDB,
32'hBE819BFE,
32'h3F0A5C7D,
32'hBEB98A8E,
32'hBE001E2E,
32'hBDF48563,
32'hBF5ECEC7,
32'h3EA719A2,
32'h3DE31120,
32'h3EDA50D6,
32'h3E0A19B7,
32'hBE00FD2F,
32'hBDAD5225,
32'h3E6EA7FD,
32'hBDA87581,
32'hBDBC8CA2,
32'hBDB44EA8,
32'h3E6BBCE4,
32'h3F8A038A,
32'h3D0E3BA3,
32'hBEEBE42D,
32'h3FA55408,
32'hBEA941DD,
32'hBEC22D47,
32'hBFC51C42,
32'hBEE98F7C,
32'h3DF7BC2A,
32'h5DE5827F,
32'h1DD6B57C,
32'h3E04AB67,
32'hBF0B88DE,
32'h3DE78730,
32'hBEE55D95,
32'h3CEE765C,
32'hBE6A1A4C,
32'h3F546520,
32'hBF4E99AA,
32'h3DC60CAD,
32'hBEC13AF7,
32'h3F1C8EF5,
32'hBEE13A16,
32'h3E4D4319,
32'hBDEBBD31,
32'h3E97D011,
32'hBE1E9850,
32'h5DE7CD10,
32'hBD834509,
32'hBE9ED27B,
32'hBE6F147B,
32'h1DED004C,
32'h3D5C2DA8,
32'h3DB8F8E5,
32'h3F4B004A,
32'hBFA8E6B7,
32'hBFD3FD83,
32'h3E3B9135,
32'hBDA3B1F5,
32'hBE06C377,
32'h3ECC7291,
32'hBE31C266,
32'hBEB10065,
32'h3CC2AFCD,
32'h3E87768E,
32'hBEB5A5D7,
32'hBFD00A45,
32'h3EEE1070,
32'hBE19E444,
32'hBF2257F9,
32'h3F38E541,
32'hBE1FE340,
32'h3ED3BBFC,
32'h3D132264,
32'hBEB56021,
32'h3D5D3A7D,
32'hBEE8DEC0,
32'hBD025A7D,
32'hBD95E588,
32'h3D6BC644,
32'hBE837C09,
32'h3E900C52,
32'h3E604AD2,
32'hBE05AA91,
32'h3ED03D00,
32'hBFA4C513,
32'hBE58997D,
32'hBF540E08,
32'hBCA1531C,
32'hBF2E4910,
32'hBEA062ED,
32'h3E64DFF9,
32'h3D69F23E,
32'hBD018F91,
32'h3E5CCCB5,
32'h3E4E402F,
32'hBFBC33C9,
32'h3DAECBE1,
32'hBF7227E2,
32'hBE96F37A,
32'h3DB18ED3,
32'hBD772D9E,
32'hBE763B26,
32'h3EC5F5BC,
32'hBEFE9F7B,
32'h3DEFFD60,
32'h3D04DB8B,
32'h5DC7905F,
32'h3C841C64,
32'h3F1622F8,
32'hBE39BC71,
32'h3E46CFF1,
32'h3EB1239F,
32'h3E4A9C8D,
32'h3DACC047,
32'hBF81EFC2,
32'hBF5EC5FC,
32'hBE691F86,
32'h3CA787EC,
32'hBFE0DC89,
32'h3DE71437,
32'hBEBB5F12,
32'hBCED3900,
32'hBE046818,
32'h3C9B84AF,
32'h3EA1FB08,
32'hBF8D99D0,
32'hBE128785,
32'hBE0E285D,
32'h3E07F434,
32'h3E3D75F2,
32'h3E5FEEFC,
32'h3D1560CA,
32'h3EABF68E,
32'hBE0E1448,
32'hBDC227A1,
32'h3E75C0AA,
32'hBD1F843D,
32'hBC913C18,
32'h3E86A448,
32'hBE79E1FC,
32'h3D169BE4,
32'h3E5E227A,
32'h3E1D1ED5,
32'hBE0F0AAB,
32'hBFA1A3EA,
32'hBFA905EA,
32'hBEFE7BF2,
32'hBE3063F2,
32'hBE3509C6,
32'h3E0988E6,
32'h175FAF92,
32'h3DE932B6,
32'hBE5C9563,
32'hBEF03FC0,
32'h3D92CB90,
32'hBF9955F2,
32'h3E15A86C,
32'h3EE665EF,
32'h3E257710,
32'h3E3F882F,
32'h3E17D83B,
32'hBD8027BA,
32'hBE4DB0A1,
32'hBE761922,
32'hBD30B9AC,
32'h3E2D95F8,
32'h075D6001,
32'hBD23C08E,
32'h3CFA5D03,
32'hBE536027,
32'h3EABB1A6,
32'h3CE45F6A,
32'h3D5202E9,
32'hBE6847E9,
32'hBE028649,
32'hBFD885CC,
32'hBE2F1279,
32'h3E113608,
32'hBE9D6571,
32'hBE5C45AD,
32'h3D658DB4,
32'h3E3156EB,
32'hBD8926A8,
32'hBD96C55C,
32'h3E54235C,
32'hBE9941FC,
32'hBD46CC8F,
32'h3E905659,
32'hBD2B1D66,
32'h3CEEEB22,
32'h3E1EE237,
32'hBDD87653,
32'h3D674E73,
32'hBE02523E,
32'h3CE124F6,
32'hBDB672C6,
32'hBD67EA15,
32'h3DA1AC32,
32'h3E009AAC,
32'h3D48438C,
32'h3E6AF2C3,
32'h3D81BC8C,
32'hBDB55D3A,
32'hBD9D0482,
32'h3CE8445B,
32'hBFCD6688,
32'hBE467771,
32'h3EB82721,
32'h3D9C796C,
32'hBE8FF953,
32'hBE284DDA,
32'h3E960301,
32'h3E384AE5,
32'h3DAA0C3D,
32'hBDC2AD11,
32'h3D453A6B,
32'hBE3670B4,
32'hBE821709,
32'h3D85DE9C,
32'h3E4FC1B4,
32'h3D6BE625,
32'hBEBD58F4,
32'h3DF427BF,
32'h3CACDF85,
32'hBEFAF0FA,
32'h3E4B58B3,
32'h3CF1A4C8,
32'hBD8087B6,
32'h3EBB29C7,
32'h3EB02BAC,
32'hBE353F94,
32'hBE5F3141,
32'hBEC2A681,
32'hBE3DCE4A,
32'h3D99DEFA,
32'hBF0195B6,
32'hBE5084E3,
32'h5DEEE8EC,
32'h3DEBCF42,
32'hBE67BFC0,
32'h0EDAE0B5,
32'h3E418731,
32'h3E01AD6B,
32'h3D2E793E,
32'hBD56DF9C,
32'hBE579311,
32'hBEB3A6E9,
32'hBE1EC2FC,
32'h3EAE37A4,
32'h3E22C126,
32'hBD7D6316,
32'hBEA44982,
32'h3D3644B9,
32'h3CD322A8,
32'hBE8B6F13,
32'hBEB9473B,
32'hBD036998,
32'hBD484056,
32'h3EB8E4C2,
32'h3E645F11,
32'hBE2E9AC6,
32'hBE64EA52,
32'h5DDECC35,
32'h3CF9588A,
32'hBEC183CF,
32'hBCF126D0,
32'hBE923C84,
32'h3DCE316D,
32'hBE887A8C,
32'h1DCCD6C7,
32'hBD33BF7B,
32'h3D212ACD,
32'h3E9504C1,
32'h3DC0A3F4,
32'hBCC23BE8,
32'hBD8A5C5B,
32'hBEF397F2,
32'hBD05FBD4,
32'hBD391AA6,
32'hBCEA1D03,
32'hBCA65B03,
32'hBDC6680B,
32'hBE3C38E4,
32'hBE38AEC2,
32'h3E241B90,
32'hBD992CB2,
32'hBD8DDBEB,
32'hBCE1E3EE,
32'h0EC8660B,
32'h3D0EF0B1,
32'hBE25C792,
32'hBD0998C5,
32'hBE8E2503,
32'h3C81F608,
32'hBECBCB87,
32'h1DDA2558,
32'hBE9D97E7,
32'hBCACDAF7,
32'h3E1A7375,
32'hBE074A43,
32'hBE824BCB,
32'hBE5E7278,
32'h3E4BCE40,
32'hBC92982A,
32'h3E36193C,
32'h3E460E98,
32'h3CD94722,
32'hBD9640E4,
32'h3E325F80,
32'h3CBA0FAD,
32'hBEE05936,
32'hBD8B45E0,
32'hBDDC3B2B,
32'hBE801A59,
32'hBEB01A83,
32'hBDDED840,
32'h3C5D8508,
32'hBD821FAB,
32'hBE91474C,
32'hBE76A563,
32'hBE204CE4,
32'hBE0C6F51,
32'hBD960FEB,
32'hBD6CB9F6,
32'hBEA49698,
32'hBE5A7FFE,
32'hBEE6658C,
32'hBD0B1145,
32'h3E444761,
32'h3D277901,
32'hBCCB544E,
32'h3D8179E1,
32'h3E3A9F69,
32'hBCA76002,
32'hBECE0292,
32'hBD402F88,
32'h3E65E2B4,
32'h3E20EE25,
32'h3DEE93A9,
32'h3D861F5F,
32'hBFDBC430,
32'hBD10D461,
32'hBDB3B5F0,
32'hBEB2E122,
32'hBD8FB765,
32'hBE29438E,
32'h3CA7D3D5,
32'h3C97D383,
32'hBEB2DAFE,
32'hBEF325F5,
32'hBEC7EAAD,
32'hBE3FD12E,
32'h3EEDD08B,
32'hBE0EBC72,
32'hBE9A9F8F,
32'hBE344AE6,
32'hBE84B6C6,
32'hBD3555A7,
32'hBD870F11,
32'h1753E19B,
32'hBE4ED8DB,
32'hBEB10892,
32'h3DF0BE03,
32'h1DC352C2,
32'hBF8FC315,
32'h1DEA190B,
32'hBF0D1A7B,
32'h3DA2C305,
32'hBE10927E,
32'hBD7A4A48,
32'hBE14ACCD,
32'hBE07F166,
32'h3D531C08,
32'hBCB6774B,
32'hBE9CA4AA,
32'h3C8859BB,
32'h3D599BC2,
32'hBC5AEE6E,
32'hBF09136D,
32'hBF0262A8,
32'h3D70DE26,
32'hBE3442D5,
32'h3E8810F9,
32'hBC9C35CB,
32'hBE72C49E,
32'hBE2E87D6,
32'hBE00C1DD,
32'hBE2EDE4E,
32'h3E291DC0,
32'hBE1087FF,
32'h3DC9690D,
32'h3E580DA0,
32'h3D790F24,
32'hBE33CBC3,
32'hBF283D22,
32'h3E8078DB,
32'h3E662E28,
32'h3CF296BA,
32'hBEAD6335,
32'hBC2309A4,
32'hBE9C2C31,
32'h3D136654,
32'h3DB7C4E4,
32'hBDB8AC23,
32'hBF5BD6F9,
32'h3DFAC799,
32'hBD5F8E9D,
32'hBDF99D64,
32'hBD5C52A4,
32'hBEEC7787,
32'h3E0725A0,
32'hBE4C2E05,
32'h3ED411EF,
32'hBE4F5D56,
32'hBE80216F,
32'hBED7B649,
32'h3ED3F576,
32'h3C93DB94,
32'h3DF46A0B,
32'h1DFA987D,
32'h3E21A970,
32'hBCA647AB,
32'hBD278791,
32'hBE31BCE0,
32'hBF240AB1,
32'h3E6510D6,
32'hBEFDF283,
32'h3E9B1928,
32'hBC25BCC0,
32'h3E4D1F8B,
32'hBEA6EACF,
32'h3DB6A7CF,
32'hBE1DC135,
32'h3E94BFFB,
32'hBF5D1F20,
32'hBEA1427B,
32'hBD3866FB,
32'hBCF419EF,
32'hBD954338,
32'hBDB5E774,
32'h3EE291F4,
32'hBE50DD5D,
32'h3ECF7667,
32'hBE1FCF2C,
32'hBE656E5D,
32'hBE3799A8,
32'hBDEA4DF6,
32'h3DA664F1,
32'h3D2C8A57,
32'h3DDB5406,
32'h3DBE18FA,
32'h3E11F235,
32'h3D8FA91E,
32'hBD8248DF,
32'hBF50E4AE,
32'hBE26E429,
32'hBF7FC064,
32'h3E8F0041,
32'hBD2A01A2,
32'h3E89F70C,
32'h3F2C425B,
32'h3E822FDB,
32'h3DD6BB70,
32'hBE312943,
32'hBEB6AEE9,
32'h3EFCA876,
32'hBD6CD52E,
32'hBDAA82F6,
32'hBD1CE279,
32'hBE1FCE30,
32'h3EC68172,
32'hBD52142E,
32'h3F472858,
32'hBED7816F,
32'hBE806551,
32'hBE013659,
32'hBE24F9D6,
32'hBDEBCCF1,
32'hBEEF1D67,
32'hBE096F1B,
32'hBED52CA1,
32'hBEB9AE20,
32'h3E56F2CD,
32'h3E06EFE4,
32'hBEB05A33,
32'hBD9EB183,
32'hBE170434,
32'h3E9AAB3D,
32'h3EEF4D4A,
32'hBD4A966F,
32'h3E69C71B,
32'h3E3C4C58,
32'h3E63EA6C,
32'hBED5CDF3,
32'hBFAB6BBF,
32'hBE05BCC7,
32'h3CD7A759,
32'h3D01A950,
32'hBF0D29FC,
32'h3D95A372,
32'h3E1D14F9,
32'hBD9CB103,
32'h3EFDA91D,
32'hBD8DECED,
32'hBDCA0E82,
32'hBE18C395,
32'h3F07AA3A,
32'hBEFC48BB,
32'hBED8EE76,
32'hBE10D321,
32'h3E825A49,
32'hBF3CAB3E,
32'h3DDFBCA2,
32'hBE27292F,
32'hBE4CD722,
32'h3DF3A652,
32'hBEE60996,
32'h3E248E47,
32'hBC4B55F2,
32'h3EA78F7C,
32'h3F099BAD,
32'h3E89391C,
32'h3D34E47F,
32'hBE32E48B,
32'hBF7B4D3E,
32'hBD605747,
32'h3CA0F740,
32'hBC4B3006,
32'hBE43DA72,
32'h3DF2C7F2,
32'hBE040ED1,
32'h3DC32D97,
32'hBEB97D33,
32'hBE851EF2,
32'hBE553372,
32'hBE6B5333,
32'h3EADC5DA,
32'hBD5B56AC,
32'h3E443698,
32'hBE216DC5,
32'h3DA0BD05,
32'hBEDFBF4A,
32'h3E59A3CE,
32'h3E2C8EF1,
32'hBF05F2B0,
32'hBF0F1D53,
32'hBDB9A6FA,
32'hBD77C0FE,
32'h3EC82ECA,
32'hBE87B23E,
32'h3EB76777,
32'hBCBEAD97,
32'hBEA9786F,
32'hBF817FB9,
32'hBF617EE9,
32'h3E339556,
32'h3D66D93D,
32'h3CA69583,
32'hBE2CED5F,
32'h3E408558,
32'h3EC1F135,
32'h3C0FA3EF,
32'h3D4EEA8E,
32'hBDEB4BFF,
32'hBEE1899F,
32'h3CFEB765,
32'h3DB5B05C,
32'hBD4DA513,
32'hBF2EA57D,
32'h3E85368C,
32'hBE82BFDA,
32'hBE7F36DC,
32'hBD9E47D8,
32'h3E20620C,
32'hBF25208D,
32'hBDA3ABF7,
32'h3EBE653A,
32'hBE94440F,
32'h3E794D5A,
32'h3D51712C,
32'h3D80AE1C,
32'hBF124D28,
32'h3CB6A954,
32'hBF84ED19,
32'hBF57B0C6,
32'h3D37E57D,
32'h1DD2FE00,
32'h3D10C01D,
32'hBD923BE4,
32'h3ED2F8D8,
32'h3E04D951,
32'hBE7CD7D3,
32'h3E9034AB,
32'h3DCE01E0,
32'hBE500FAB,
32'h3E462F8F,
32'hBE774D99,
32'h3E051392,
32'hBE6B6A83,
32'hBEF6CCE0,
32'h0ED10177,
32'hBEF8D83E,
32'h3EF5275C,
32'h3E44E12F,
32'hBDC6EFFC,
32'hBDAABCA2,
32'h3EDF40ED,
32'h3D138C9B,
32'h3E2E24D3,
32'hBF156D93,
32'h3EB7DFC2,
32'hBE9802D3,
32'h3F57672B,
32'h3EDB6B4A,
32'h3DB40FC3,
32'h3F01918E,
32'h3D1A8AE1,
32'h3C19CDEC,
32'hBF89B554,
32'hBDCB5B8F,
32'hBD54A02E,
32'hBD000B2C,
32'hBEDFF578,
32'hBF3C47AA,
32'hBD8A312D,
32'h3D051219,
32'hBF70D8BE,
32'h3E6508EC,
32'hBE3AF2AA,
32'hBE7B50C6,
32'h3E8A739F,
32'hBF538B08,
32'h3F81B647,
32'h3DF5E478,
32'hBDAF72E7,
32'hBF97CF58,
32'h3EE93621,
32'hBCD1BC67,
32'h3E564700,
32'hBF5FB237,
32'hBDEF873E,
32'hBF086945,
32'hBE8652FB,
32'hBF2FF727,
32'hBD6E3AC5,
32'h3F44E2F5,
32'h3D669358,
32'hBC80D60D,
32'hBF483338,
32'h3EE6226B,
32'h3EF40F4D,
32'h3DF32F39,
32'h3F67B6E6,
32'hBE9FB400,
32'h3DAF6061,
32'hBE10900E,
32'hBF4502C1,
32'h3E30C5C0,
32'hBF4FC072,
32'h3F5419E4,
32'hBE2B9CF1,
32'hBC3E8E14,
32'h3EFC4DD1,
32'hBEC1E526,
32'h3EC5FB86,
32'hBEB20FBB,
32'h3CF19EEE,
32'hBD4595D3,
32'h3F48BF12,
32'h3E1083B8,
32'hBE390805,
32'hBE00BA9B,
32'hBDE27C8B,
32'hBE73D5E4,
32'h3F08F26F,
32'h3FA333BD,
32'hBD9B3EBE,
32'h3D90C628,
32'h3F3C922D,
32'hBF06CAC9,
32'h3ECB7E58,
32'hBE776E58,
32'h3FCB7CE5,
32'h3E0583EB,
32'h1CD518A,
32'hBE4F8D69,
32'hBF11280E,
32'h3C9EB105,
32'hBF27F825,
32'h3F691AD3,
32'hBD86D1B0,
32'h3EC52E78,
32'h3E57D45A,
32'hBF3C13F6,
32'h3F2BEDFA,
32'hBEB6D1BD,
32'h3F542FF5,
32'h3DDEA3CC,
32'h3DEDE7E3,
32'h3FEC2DAC,
32'h3D492A09,
32'h3E5C67E6,
32'hBEFF0D25,
32'h3D8ABCFA,
32'hBD810A01,
32'h3F79A387,
32'h3D1496B0,
32'hBDA92022,
32'h3FB3C61F,
32'hBFA2219E,
32'h3C106724,
32'hBF7C2EFB,
32'h3EACD3B7,
32'h3F4A9F6C,
32'hBF9661AD,
32'h3ED231BC,
32'h3F26BC22,
32'h3ED33156,
32'hBE256E23,
32'h3F5D2B01,
32'h3E45CF2F,
32'h3D8D92ED,
32'hBF2CFE8A,
32'h3D932D23,
32'hBF2409D6,
32'h3F67F8E8,
32'h1DDCFE69,
32'h5DEC5662,
32'h3C285D52,
32'hBD27856A,
32'hBC9BBDA2,
32'h5DFF1A27,
32'h3DA1F267,
32'h3C89E1E6,
32'hBDBA136C,
32'hBCDB7294,
32'h3DAE56E1,
32'hBD31BE11,
32'h3DC312D9,
32'h3CF666D8,
32'hBD6D5C6A,
32'hBD848165,
32'h3D156F39,
32'h3CDF2FEB,
32'h3D4AAC9E,
32'h3DDD9884,
32'h3CEFB4A3,
32'hBDF7F5D0,
32'h5DC37EAB,
32'hBD9A64CA,
32'h3D6E0A15,
32'h3CCF1E12,
32'h3CDD0BA3,
32'h3D8A546C,
32'hBD08E9B1,
32'hBCC5E574,
32'h3CEB36A5,
32'h3D8E6712,
32'hBD964715,
32'h3D4EF308,
32'hBD461C13,
32'h3D99552F,
32'h3CAB0FB9,
32'hBD4593EA,
32'h3DBB548E,
32'hBD68177C,
32'h3D9A0801,
32'h1DE8894B,
32'hBC984228,
32'hBD040978,
32'h3C4C0CEE,
32'hBC016708,
32'hBCD4D164,
32'h3D043564,
32'h3CAA09D4,
32'hBD3D7822,
32'h3CBB0A76,
32'h3CF7E207,
32'h3D849CC5,
32'h3C8B3F78,
32'hBD8CF870,
32'hBDB48D14,
32'h1DC20642,
32'h3C2497AA,
32'h3D7E06FC,
32'hBDEA4FAA,
32'h3C8AF14B,
32'h3CA08B72,
32'hBC8B70CA,
32'hBD4255C7,
32'hBD587600,
32'hBD2F2A71,
32'hBDC5A209,
32'hBD3EEABF,
32'h3CEE9444,
32'hBDDECC6B,
32'h3D44A876,
32'h3CB7F00B,
32'h1757156B,
32'hBD90AD03,
32'h1DEDFFF8,
32'h3CB5D621,
32'h3CB5EC5C,
32'h3D456DC8,
32'h3D91D1D7,
32'hBD81B704,
32'hBD8B3D1F,
32'hBD16B9F6,
32'h2ED2FD6C,
32'hBD7C1F11,
32'h3C42D0FB,
32'hBCF22D00,
32'h3D62578F,
32'hBD34D5C1,
32'h3CA5818F,
32'h3D48CCFF,
32'hBE145229,
32'h3EC968E1,
32'h3F202BCF,
32'hBE0835E3,
32'hBEC14C7F,
32'hBE864568,
32'h3EB9E0D9,
32'hBEE03BFD,
32'h3E3C5739,
32'hBD32BE96,
32'h3D81B6C0,
32'hBD051992,
32'hBECB0567,
32'h3F1C8A62,
32'h3EB2F527,
32'hBE4C5E4B,
32'h1DE4B2A8,
32'h3D40F380,
32'h3C845911,
32'hBD30DF02,
32'hBE7195CA,
32'h3CA58D68,
32'hBDC8D1FE,
32'hBF0262CA,
32'h3EE3DE12,
32'hBDD02196,
32'h3F3415BB,
32'h3F3D1FFF,
32'hBEA81C51,
32'hBE665CAE,
32'hBF7BC210,
32'h3EB208DC,
32'hBEAB3552,
32'hBF4868B6,
32'hBE879A95,
32'hBF55A2D6,
32'h3EE7C449,
32'hBE8E437E,
32'hBE8EF276,
32'hBC7B3D09,
32'h3D71A17D,
32'hBDDB5B0D,
32'hBF5113DD,
32'hBF207469,
32'hBE7FE2D5,
32'hBE827489,
32'h3F9ECD05,
32'hBF373DB1,
32'h3C954E6E,
32'hBED7B271,
32'hBF0E857E,
32'h3E8E6535,
32'hBDC1DC9E,
32'h3E2942D7,
32'hBEA23436,
32'hBF54FDED,
32'h3ED0C039,
32'hBD7B86A0,
32'h3EB78DA2,
32'h3E7F40E5,
32'h3E2FCCF7,
32'h3F0DD08E,
32'hBF04748F,
32'hBF96A79F,
32'hBD65BBA8,
32'hBF19F690,
32'h3E8DFED2,
32'h3E50888D,
32'hBD825F74,
32'hBF36BEFB,
32'h2EDEAC76,
32'hBC86ABB9,
32'hBF506D57,
32'hBE33E8A5,
32'hBE35B0FC,
32'hBD160805,
32'h3E2143E9,
32'hBF453AAD,
32'hBFA738D0,
32'hBF886484,
32'hBFA85C57,
32'h3F252679,
32'hBCBF8A94,
32'h3EF88EB4,
32'h3F14F4AD,
32'hBD8FAC9F,
32'h3F47A68B,
32'h3F444CB4,
32'h3CC5B2AA,
32'hBE92AA96,
32'h3F0EB12E,
32'h3ED4359E,
32'h3DED828F,
32'h3ED1345E,
32'hBE299B49,
32'h3F1E8DD8,
32'h3E803E9D,
32'h3D2D49B6,
32'h3D8A2697,
32'hBF717E12,
32'hBD2886CB,
32'hBCF70D02,
32'hBDBB3221,
32'h3EB800C9,
32'h3EAA776E,
32'hBDC3C52B,
32'h3D806789,
32'hBF13CB8F,
32'hBF2563B8,
32'hBF038CC0,
32'hBF490745,
32'hBDDE477C,
32'hBEADDE05,
32'hBEE7728A,
32'h3F3128B8,
32'h3F805DA3,
32'h3F59639E,
32'h3EFFDAAE,
32'h2EC59695,
32'hBEE83031,
32'h3E61A45F,
32'h3EF8B256,
32'h3EF5ECE2,
32'h3E6D6504,
32'h3EC2FAC2,
32'h3E4940AE,
32'h3E61A6AA,
32'hBEC661D2,
32'hBDCD3E56,
32'hBDF3F895,
32'hBCD8F2AE,
32'h3C73A75D,
32'hBE1A3D5A,
32'hBE5D8BD5,
32'h3E975B07,
32'hBD92C3F3,
32'hBE32CFD6,
32'hBE972C52,
32'hBEBCC4CE,
32'hBF07208D,
32'hBCFB4B20,
32'h3C9DFA2F,
32'hBF394DC8,
32'hBD1E7CE9,
32'h3E8FF08A,
32'h3F702DD9,
32'h3F039273,
32'h1DF09C85,
32'hBC55DD92,
32'hBF5FC4AF,
32'hBE8D497B,
32'h3EDEDBF7,
32'h3EFC4277,
32'h3DA767B8,
32'h3F2B2848,
32'h3DD8A593,
32'h3DD05F72,
32'h3CC49722,
32'hBEAC1F6B,
32'hBF4D924B,
32'h5DE932C7,
32'hBDAC8A82,
32'h3EB620BC,
32'h3D3AD6EC,
32'h3E813BB8,
32'hBDB4AD93,
32'hBE391DD8,
32'hBC42E663,
32'hBEB23D9B,
32'hBF5D3647,
32'hBEC3DCB0,
32'h3E4C3BA5,
32'hBFAF4FF4,
32'hBC4A1A21,
32'h3D4F0E28,
32'h3F365A1E,
32'h3EC972F9,
32'h5DDD7D16,
32'hBEABC933,
32'hBE18B545,
32'h3E8F0937,
32'h3DED2781,
32'h3E1EF71D,
32'h3E5F9A65,
32'hBD6C28DE,
32'hBD5ED606,
32'h1750E129,
32'h3E359EEF,
32'h2ED5185A,
32'hBD6A8602,
32'hBCF4210D,
32'hBD4962B8,
32'hBD0B05F3,
32'hBE871A6F,
32'h3E1C5576,
32'h3D4415D0,
32'h3E2FB35A,
32'hBD2B1E1D,
32'h3D84DF9B,
32'hBF23DE49,
32'hBEFE3120,
32'h3D8EE592,
32'hBF784FF8,
32'h3C9173F6,
32'h3CD0C123,
32'hBEA505EF,
32'h3DD8916B,
32'hBE8E1513,
32'hBE9F67A4,
32'hBF17BC94,
32'hBE10C274,
32'hBC256AF4,
32'h3ED296B1,
32'h3E2F3C3B,
32'hBE0BCCBC,
32'h3E94DE46,
32'h3EB424DC,
32'hBDC6DD0C,
32'hBE06DD67,
32'hBE1223DC,
32'hBDCADBCA,
32'hBC199FA2,
32'hBDEEFBA6,
32'hBD8CEBCC,
32'h5DE63E87,
32'hBDECF6FE,
32'hBDD0FEC0,
32'hBE58AD40,
32'hBDAA531B,
32'hBD8378C6,
32'h3A11F83,
32'hBD592BA0,
32'hBE9A0E5F,
32'hBE805520,
32'h3DEBA32A,
32'hBD7E4EB0,
32'h3E9B6435,
32'h3E36E16C,
32'hBF59F20F,
32'hBF23D87E,
32'h3C1CFF63,
32'hBDD7D883,
32'h3E49ED81,
32'h3EDE03D0,
32'hBE53DE12,
32'h3E0DB1F4,
32'h3E2187C4,
32'h3E348ECD,
32'hBF04D1FA,
32'hBE645529,
32'hBD0B78EB,
32'hBD94B390,
32'h3E64470B,
32'hBD3D2728,
32'hBE2E8278,
32'hBEBE267F,
32'h5DEABE89,
32'hBE42E610,
32'hBC4C790C,
32'hBDA97652,
32'hBCA09E74,
32'h3CF04FED,
32'hBF40769A,
32'hBF0B3442,
32'hBE23F478,
32'hBCB8481D,
32'h3DE1EB11,
32'h3E90F8DD,
32'hBF818689,
32'hBE843F19,
32'h3E673548,
32'hBEB4968F,
32'hBD5FA6E5,
32'h3DCFE8DF,
32'h3D4A8AA6,
32'h3D94A2D3,
32'h3E04AF46,
32'hBDAC3F72,
32'hBECC467D,
32'hBE021DD3,
32'hBD275E13,
32'h3C2F2BC5,
32'hBDD9B9C6,
32'hBE8019C2,
32'h3E02050C,
32'hBE5D9E06,
32'hBE5CD9EF,
32'hBDA46525,
32'hBE206FBC,
32'h3EC5B957,
32'hBD0A6CAC,
32'h3E62DC08,
32'hBF3FBCEF,
32'hBEE3A9FB,
32'hBD948EA3,
32'hBE08806D,
32'h3E8D0B7D,
32'h3E63E30F,
32'hBF713DFA,
32'hBE74F248,
32'hBD34049D,
32'h3CFBB009,
32'hBCBD72B5,
32'h3C86F706,
32'h3E19FC99,
32'h3D58CD88,
32'h3D027DDA,
32'hBC60BF0A,
32'hBEE80C86,
32'h3DF1FFA1,
32'hBC30B471,
32'h3CBBD603,
32'hBF0BFF11,
32'hBEE25BAF,
32'h3DBACDF4,
32'h3D6E8871,
32'hBE3F55CA,
32'h3D2CBFC1,
32'hBE535DEA,
32'h3C740AB5,
32'h3C177FDB,
32'h3CD858F5,
32'hBD4822D1,
32'hBDCFD972,
32'hBE294CD1,
32'hBE8263F8,
32'h3DB1C01D,
32'h3D152B61,
32'hBEFDCC7F,
32'hBEE0EFA9,
32'h3EB8CF45,
32'h3E61E246,
32'h3D936793,
32'h3D0C807D,
32'hBE3762BD,
32'hBE4FCDF1,
32'hBD8873C5,
32'hBDCF1C94,
32'hBEAB3DC2,
32'h3D824AC5,
32'hBD4DF357,
32'hBDBE6CD9,
32'hBF22A285,
32'hBED3AAB6,
32'hBE2A8401,
32'h3D8A177F,
32'hBF08F654,
32'hBDB5525E,
32'hBE2560F4,
32'hBEEB41CD,
32'hBE693C81,
32'hBDF0AFE9,
32'hBF251F32,
32'hBE1B9DC8,
32'hBC38BA38,
32'h3D8A820D,
32'h3E211058,
32'hBCF8E139,
32'hBF59222B,
32'hBEDBDF7E,
32'h3D3B4208,
32'h3C3CF6E6,
32'h3DD97FAD,
32'h3E8FF64D,
32'hBFCEC6C8,
32'h3CEEC108,
32'h3D5250C7,
32'hBE643A9D,
32'hBDCE8C1C,
32'hBE3A72AF,
32'h3D0E2D68,
32'hBCAE3432,
32'hBEB074EE,
32'hBEAA3B38,
32'hBE89962E,
32'hBE5D029A,
32'hBE8FB55A,
32'h3D951E34,
32'hBE7D4096,
32'hBE88AC88,
32'hBE4F4A03,
32'hBDFFDD32,
32'hBF4B675F,
32'hBD864FD4,
32'hBC729735,
32'hBE024895,
32'hBCDBA17D,
32'h3D0565F5,
32'hBF947F39,
32'hBE99AA4B,
32'hBE1A6D91,
32'h3EA7DA73,
32'h3D926CA5,
32'hBD917BFA,
32'hBF1D4CFA,
32'hBCF74B11,
32'h3E61DE12,
32'h3E3A19EE,
32'hBE826002,
32'h3E71C12B,
32'hBDEF5357,
32'hBD0F8872,
32'hBF03FEDF,
32'hBEADDA2E,
32'h3E4D8BC0,
32'h3E264747,
32'hBD47272B,
32'hBE6A7D41,
32'hBEEBF773,
32'h3E934C54,
32'hBEB4AAD3,
32'hBE06AB6B,
32'hBF1DC338,
32'h0ED6D5FF,
32'hBE262503,
32'hBC02DD91,
32'h3E42B4AD,
32'h3D896F42,
32'hBF1B3EE2,
32'hBDBCE0DD,
32'h3EDE5407,
32'h3E82A475,
32'hBEC58327,
32'hBDB0EF54,
32'hBFA991A1,
32'hBD93D391,
32'h3D88E29E,
32'hBD7A7090,
32'hBEA29238,
32'h3E5D6DE3,
32'hBD569ADA,
32'hBDE85E08,
32'hBFA9F73F,
32'hBF00FF6E,
32'h3C813C66,
32'h17555957,
32'h3EAA0753,
32'h3D21AC3F,
32'hBED44156,
32'hBE9F1B5B,
32'h3EC77FCF,
32'h3CC672AC,
32'hBF042FBA,
32'hBE8A753B,
32'h3E2FE389,
32'hBE2AB24B,
32'h3D0E1141,
32'hBCE60645,
32'hBF2398EA,
32'hBE25D47E,
32'hBEAF76DF,
32'h3EFF8451,
32'hBEB75C30,
32'h5DC3BCA8,
32'hBFE71063,
32'h3E7AA8D5,
32'hBED402DC,
32'hBE9FAA1A,
32'hBEFCCBD2,
32'h3E17239E,
32'hBCA9A567,
32'h5DE601C9,
32'hBF5AE729,
32'hBE0AE140,
32'h3EB82FED,
32'h1DF0F5DA,
32'h1DC74EAE,
32'hBE3F2A5E,
32'hBE882B03,
32'hBD6735AA,
32'h3E7EAF2B,
32'hBC9B573A,
32'hBF3CA028,
32'hBCF3AB8A,
32'hBE450827,
32'hBE851E6F,
32'h3DA0017B,
32'hBECF9E6A,
32'hBF842A68,
32'hBC4FC3CA,
32'hBEC559D1,
32'hBD3C5B0D,
32'h3EBAB925,
32'hBE4C49F8,
32'hBF0BAE2E,
32'h3E93C6D0,
32'hBE18B34B,
32'hBEF9ECE1,
32'hBE885CD9,
32'h3E767B55,
32'hBC819DF0,
32'h3D784A68,
32'hBF4DC7E5,
32'hBEACE7B7,
32'h3E868BF6,
32'h3C3A8BE4,
32'h3E0B20CC,
32'h3DA5780A,
32'hBE732156,
32'h3E9850A8,
32'h3EA78F36,
32'hBF074C2D,
32'hBEC0DAEC,
32'hBE2C6DAB,
32'hBCB2F9B7,
32'h3DAB0A57,
32'hBE2DDE60,
32'hBC889F39,
32'hBE907ABE,
32'h3ED4D02F,
32'h3D8B636D,
32'h1DE30272,
32'h3E285035,
32'hBF7BDB59,
32'h3DB3306F,
32'h1DE9E205,
32'h3E8A2048,
32'hBF3A1FA9,
32'hBFA4B4F0,
32'hBEE71CFD,
32'h3CA5E8F9,
32'hBC99C49F,
32'hBF5DC1E9,
32'hBE5FD504,
32'h3ED69061,
32'h3DC4FF54,
32'h3E82743C,
32'hBE664080,
32'hBE57ACCF,
32'h3EA1C8E0,
32'hBE360751,
32'hBE864B9C,
32'hBD1646D5,
32'h1DD0EC01,
32'hBCC2762B,
32'hBF8F1D0F,
32'hBE03F667,
32'h3E6A99ED,
32'hBE340B2F,
32'hBDC8A47F,
32'hBEFD107E,
32'h3E8876B6,
32'hBE76253A,
32'hBF5CA29A,
32'h3EB7743A,
32'h3EBD97B9,
32'h3DB94022,
32'hBF949C64,
32'hBEEAAD36,
32'h3DDF869D,
32'h5CD8144,
32'hBDCB3B34,
32'hBF6667A4,
32'h3E040080,
32'h3C19A76F,
32'h3E1CF761,
32'h3D7A0F87,
32'hBE9BEE40,
32'hBEB791DC,
32'hBDF2DEB5,
32'hBED81F6B,
32'h3D268380,
32'hBE9A6B28,
32'hBECA5837,
32'hBCCBB7CA,
32'hBF03A41A,
32'h3E8AB770,
32'h3E68DBC8,
32'hBF68A1F3,
32'h3F150F44,
32'hBE0DAB76,
32'hBE05B59D,
32'hBD52526F,
32'hBF58D5EC,
32'h3DEC4D20,
32'hBEA511B4,
32'h0EDE543A,
32'hBFC72B30,
32'hBE4317A4,
32'hBF017341,
32'hBD10E105,
32'h3D8A60C9,
32'hBF564835,
32'h3EDD3BFC,
32'h3E825586,
32'h3E2808FF,
32'h3E3E05CE,
32'h3E9EEEAA,
32'hBD81A523,
32'h3E14F517,
32'hBE76696D,
32'hBDD83896,
32'hBC849344,
32'hBEFB1445,
32'hBE8AAC42,
32'hBEF2EDD7,
32'h3E2F65B3,
32'hBE07802C,
32'hBF36CA8C,
32'h3EE12E3C,
32'h3D939FED,
32'hBEB134D8,
32'h3D5DF4AA,
32'hBEF4DF14,
32'h3D9B0B2F,
32'h3DFC8643,
32'hBEA863C6,
32'hBF8B7BE2,
32'hBF885489,
32'hBD862690,
32'h2EC02731,
32'hBCD5BA11,
32'hBF297C3D,
32'h3F4F2CE6,
32'h3EF33122,
32'h3E7C62DC,
32'h3F2B5242,
32'h3DB086C8,
32'hBDE12351,
32'hBF12F5EF,
32'h3F4F720C,
32'hBE05E692,
32'hBF6E6383,
32'hBEBDB129,
32'h3E62C194,
32'h3E050DFE,
32'h3F45ADDD,
32'hBDB01816,
32'h2EC94C5E,
32'hBF0FEF5A,
32'h3DCEB7CF,
32'hBF900895,
32'h3F18710C,
32'hBFBFFA84,
32'hBD6ABEE7,
32'hBE99DF35,
32'hBE020616,
32'hBF1B789D,
32'hBEF6D490,
32'hBE03CAF6,
32'hBD9A9CC6,
32'h3D497B40,
32'hBF301676,
32'hBE0A21ED,
32'h3F1A1829,
32'h3E1127C4,
32'hBF1D9DDE,
32'hBE60972E,
32'hBE425AD5,
32'h3D910EE6,
32'h3F5786D7,
32'h3E1B6A29,
32'hBF07119B,
32'h3D8C5425,
32'h3CFBDEBE,
32'hBF3500FF,
32'h3ECEFB4C,
32'h3D71DEB6,
32'hBF2A8DD8,
32'hBF20EA1F,
32'h3F004C4C,
32'hBDA82549,
32'h3F117CDB,
32'h3E86CABC,
32'h3F0A8BDC,
32'hBF901E82,
32'hBF28DEFE,
32'hBEA9B3F5,
32'h3D2432C3,
32'hBE163D63,
32'hBC2FA703,
32'hBCB0D8A3,
32'hBEE87C3E,
32'hBEC46B43,
32'h3F02ACC7,
32'h3F89A3A3,
32'h3FA6EEFF,
32'hBEB06565,
32'hBF1C9424,
32'h3C1EF372,
32'h3E773F73,
32'h2ED8E652,
32'hBE072C71,
32'h3F3090B4,
32'hBF1E191C,
32'h3F966E5B,
32'h3EB97BB2,
32'hBD6E7A8F,
32'hBF3C91EF,
32'h3DE24CB6,
32'h3EA5D9F9,
32'hBD9AAC55,
32'h3D160050,
32'h3F249D8A,
32'h3DDDC9CA,
32'hBEF682B0,
32'hBF26198C,
32'hBE76DA1E,
32'hBE283501,
32'h3DD6FE70,
32'h1DFFDB85,
32'h3A32584,
32'h3F1C90C1,
32'hBFB25B3F,
32'h3D2AAAA0,
32'h3F97B821,
32'h3F6702F8,
32'h3F4E8011,
32'h3EA609B0,
32'h3EC9C49E,
32'h3F7D14E3,
32'hBF1C5993,
32'hBDA24D14,
32'h3F8B7A6C,
32'hBF105151,
32'h3F04A5B3,
32'hBE107634,
32'h3EB06692,
32'hBEF02B91,
32'h3EEA43D6,
32'h3F8A9734,
32'h3D1A052C,
32'hBEA527D3,
32'h3EFC75CD,
32'h3E2B50AC,
32'h3E8DA1F3,
32'hBE11115C,
32'hBE58A63C,
32'hBE9ED76F,
32'h3F8A1525,
32'hBD3440D9,
32'h3D52BE60,
32'h3F716812,
32'hBFC10704,
32'hBE6CA7E3,
32'h3E4BAE87,
32'h3ED99423,
32'h3F59FBA4,
32'hBEAC6FBD,
32'h3F448D9F,
32'h3F1D3B2C,
32'hBF2411CE,
32'hBCD47047,
32'h3D50255C,
32'hBD49673A,
32'hBC5DE722,
32'hBF31E51B,
32'h3CE141A1,
32'hBF308E4C,
32'h3F587F2F,
32'h1753EFA5,
32'h3D291AC3,
32'hBC95C2B7,
32'hBD8AC442,
32'h3D2739E0,
32'hBDB41A35,
32'hBD45617E,
32'h3D4FC70A,
32'hBD3FEE90,
32'hBDDD68EB,
32'h3D80296C,
32'h3DD0C93F,
32'h3D18A80C,
32'h3D8FFE8D,
32'h3CC44792,
32'hBCE4EAAF,
32'h3D506387,
32'h3DAAB4DB,
32'h5DEE806A,
32'h3DBC948D,
32'h3C815DD3,
32'h3A38719,
32'hBCEEE2CD,
32'h3D830FBE,
32'h3D09EB10,
32'h3C68C6C5,
32'hBD847C1E,
32'h5DF14050,
32'h3DADDB17,
32'h3D8EFF71,
32'h3D0CE43A,
32'h3D38A17B,
32'hBD808FD5,
32'h3C84AA69,
32'hBD89B832,
32'hBCD3452B,
32'h3DDA342E,
32'hBD39EE17,
32'hBC8EA90D,
32'h3C51E3D9,
32'hBD63A0B9,
32'h3D81C4BA,
32'h5CCBBCD,
32'h3D5630C3,
32'h5DCB2D61,
32'hBC9F91F6,
32'hBD751B7E,
32'hBDC4CF28,
32'h3D95EF1E,
32'hBDAE6333,
32'h0EC7B059,
32'hBD309C1A,
32'hBCB48F2F,
32'hBC880E84,
32'hBC534AF1,
32'hBDB5BCA0,
32'h1DC6E4B3,
32'h5DC5C50B,
32'hBD2029B5,
32'h3DAA50E6,
32'h3CC36C74,
32'hBD1BDCDF,
32'hBCBD1CB2,
32'hBC9A1A3E,
32'h3CC559DB,
32'h2ED922B0,
32'h3CA55FF4,
32'h3C59830E,
32'h3D9B9207,
32'h3D322203,
32'h2ED6FFF8,
32'h1DDDCCF5,
32'h3DAA8B16,
32'h3CF76298,
32'h3DE6DD2E,
32'h3D1EA976,
32'h3D4F2898,
32'hBC8C3F99,
32'h3DBFA968,
32'h3DB32A98,
32'hBCCFBAE1,
32'hBC0A60C3,
32'h3DD9665D,
32'hBDC20530,
32'hBA5B2A2,
32'h3D68799E,
32'h3DDE8580,
32'hBD266E21,
32'hBD08FF11,
32'hBD775D3A,
32'hBC167AC8,
32'h3DA13FC3,
32'h3EC6A35A,
32'h3C0DE8FA,
32'h3E46DBBD,
32'hBE9CF30D,
32'h3EB596E3,
32'h3DB180C7,
32'h3C6928C7,
32'h3CB12FC1,
32'hBCE7E1F4,
32'h3D464368,
32'h3D581E6F,
32'h3E3A9893,
32'hBE0E2863,
32'hBE0106BC,
32'hBD6DE5B8,
32'h3D353A17,
32'hBDADF984,
32'hBD7D6A04,
32'hBDF177C2,
32'hBE5E3AF2,
32'hBD4C1FB1,
32'hBE90D146,
32'hBD3C1E9A,
32'hBDFD9884,
32'h3E548F76,
32'hBC90F513,
32'hBE3C6C64,
32'hBE76A69A,
32'hBEF94B73,
32'hBE0E6839,
32'hBEB0FB95,
32'h3DCDCEBA,
32'hBEC1464D,
32'hBE3114D7,
32'h3E9479B1,
32'hBEB137ED,
32'hBF24740D,
32'hBC5042D7,
32'hBC0F5056,
32'hBCA123F2,
32'hBEA5EAA8,
32'hBFABDF46,
32'hBDAE8EEE,
32'hBF89AE26,
32'hBE895317,
32'h3CBF3300,
32'hBF2ECD74,
32'hBCAE8AD0,
32'hBE48C2D9,
32'h3EA189AB,
32'hBE43DE23,
32'hBEDA18CD,
32'h3F257233,
32'h3D3CE042,
32'h3F7C90F7,
32'h3C2103BC,
32'h3E6CADAA,
32'hBCDF7C7F,
32'hBE19ACB4,
32'hBEA58047,
32'hBED29A21,
32'h3EF7F54D,
32'h3EED8696,
32'h3F768D3A,
32'h3DB9AF98,
32'hBDE7A5E0,
32'hBF465678,
32'h3D3DE5F4,
32'h2EC88DFD,
32'h3D7FCCA9,
32'hBF70A38E,
32'hBF8D0F94,
32'h3E36EAD5,
32'hBEDFCB57,
32'hBF0BAC7E,
32'hBEC44EFE,
32'hC00278EF,
32'hBEA0F0C4,
32'hBEF4D67D,
32'h3F1A1547,
32'hBCC60B9E,
32'hBF1058BA,
32'h3F554443,
32'h3F5AD0FB,
32'h3ED2375A,
32'hBE3FF92C,
32'hBD07FD6C,
32'h3D56A2C9,
32'h3ECA7B6A,
32'h3E819657,
32'hBEA47DF5,
32'h3F68699C,
32'h3EB7BD57,
32'h3F4F3A39,
32'hBDCAEB4A,
32'h3DA0DF2F,
32'hBF9344EA,
32'hBE9994A2,
32'h3DBCBEED,
32'hBDD1843F,
32'hBF70A671,
32'hBF789B7F,
32'h3E84A07A,
32'hBD03A3A0,
32'hBEE204BB,
32'h3E4A4372,
32'hBF15AE47,
32'h3DB7ED44,
32'hBEC5CDDD,
32'h3F1A444E,
32'hBD2BE0B4,
32'hBF056628,
32'h3EC66CFE,
32'h3F691848,
32'h3EC48E59,
32'h3ED97C00,
32'hBF346BC7,
32'h3F02D780,
32'hBD3BC3B3,
32'h3E01BE77,
32'hBE938CC4,
32'h3EF13F44,
32'h3F0BD16E,
32'h3D12A2CE,
32'h3E43ECDB,
32'hBE870886,
32'hBF1C71E2,
32'h3F55A1C7,
32'hBC3A2541,
32'h3D923539,
32'hBFAFE7ED,
32'hBFC87BF8,
32'hBE2A564D,
32'hBC0C8FB7,
32'hBF4472B7,
32'h3F3ACE22,
32'hBF77F847,
32'hBD3B7D20,
32'h3DCF7746,
32'h3EEB2E18,
32'h3DBEBDB5,
32'h3EA48E59,
32'h3EAB33E6,
32'hBD59293B,
32'h3CE1BF6D,
32'hBDC06833,
32'hBF57B942,
32'hBF364119,
32'hBF021E6D,
32'h3ED22BBB,
32'hBE58E199,
32'h3DA57923,
32'h3F17EEAF,
32'hBDCEBF44,
32'h3D222907,
32'h3D77D756,
32'hBEFB827B,
32'hBF12552C,
32'h3D3C2BE8,
32'hBC1FB80F,
32'hBFA6967F,
32'hBF54F886,
32'hBE107B26,
32'hBE601D49,
32'hBF3F4CF6,
32'h3ED21E17,
32'h3DE3997E,
32'hBF6FFF95,
32'hBEE41339,
32'h3EEF6628,
32'h3DB2CCBF,
32'hBE241FD9,
32'h3E55C351,
32'hBE22EAAB,
32'h3DE56FD5,
32'hBE8D2D3E,
32'hBF48426C,
32'hBF0C6A48,
32'hBEE75BF5,
32'h3E37BE2E,
32'h3E4BD0C9,
32'h0ECEC4B3,
32'h3F13DA5B,
32'hBE6545AC,
32'h3E7BD859,
32'h3E8E87BE,
32'hBEC6B0A5,
32'hBF999BDA,
32'h1DDE79B8,
32'h3C14A85E,
32'hBF763439,
32'hBF88D837,
32'hBF2FA831,
32'hBDD645DB,
32'hBF216338,
32'hBE89DEE7,
32'hBD051915,
32'hBE53B518,
32'hBEEB85BE,
32'h3E00F8A6,
32'hBE08D5C9,
32'hBD6E6787,
32'h3E26A79B,
32'h3EBFF803,
32'h3E03BCCF,
32'hBEBE891A,
32'hBF0AA5C2,
32'hBE05025B,
32'h5DE51D40,
32'hBE9586E2,
32'h3E3E9A8D,
32'h0ED34D2E,
32'hBCFD0EFE,
32'h3EA6D68C,
32'h3DEF80BD,
32'hBF43CC63,
32'hBF7A9FD2,
32'hBE0E07DB,
32'h3DBF9BD5,
32'hBD770B92,
32'hBF7E2F63,
32'hBF56FC15,
32'hBF087F96,
32'hBEEA6AB8,
32'h3EBC5C94,
32'h3EC4E703,
32'hBEC5CF70,
32'h3EA78BC8,
32'hBDA4DCF0,
32'h3CD98FB8,
32'hBFA032C3,
32'hBE81E2BB,
32'hBD1974F7,
32'h3D97D4DD,
32'h3E4D17A9,
32'h3E2ACFAB,
32'hBF1AE677,
32'hBED4EB4D,
32'hBDB13A72,
32'h3DE58B37,
32'hBECF12F8,
32'h3E004BBB,
32'h3DCBBC42,
32'h3D3003D2,
32'h3EFE9534,
32'hBF1CA29A,
32'hBF61C83B,
32'hBE71ABED,
32'hBD00070B,
32'h3C14054E,
32'hBF7FDEF2,
32'hBEF4A7DD,
32'hBF055D97,
32'hBCDAC641,
32'hBE93311B,
32'hBE023423,
32'hBDEC6726,
32'h3D2502D7,
32'hBE2A99B7,
32'h3DD3DA7D,
32'hBF98D4E6,
32'h3E06EC50,
32'h3CF27E32,
32'hBCAD11A9,
32'h3D4E8A6B,
32'h3C006696,
32'hBF354458,
32'hBD5C6FAE,
32'hBDE297D3,
32'h3E5B248B,
32'hBD4E3CEC,
32'hBE6B4523,
32'h3EEF7A3B,
32'hBE615726,
32'h3E82DBA3,
32'hBF1F822A,
32'hBED8F08E,
32'hBE55F43B,
32'h3C0854AD,
32'h3D5752CD,
32'hBF423BD2,
32'hBEE931D7,
32'hBD654AD3,
32'hBD3A2152,
32'hBD2BDFFD,
32'hBE437F4A,
32'hBE116BFC,
32'h3EBD3757,
32'hBC8EFA16,
32'hBD86EB07,
32'hBFC14DF1,
32'hBC8B9C10,
32'h3E405632,
32'h3F069608,
32'h3E1B2BFF,
32'h3E7F68AE,
32'hBE023C5C,
32'hBD4A4D83,
32'h3EDDAEA4,
32'h5DD2BB6C,
32'h3E0F36EC,
32'h3EAD5BD3,
32'h3F386237,
32'hBD1C9FEE,
32'hBE83EBAE,
32'hBF3277DE,
32'hBDEF1F0E,
32'hBE926B84,
32'hBD3B2000,
32'h3C0030CC,
32'hBE90E9A7,
32'hBF43575A,
32'h3D3D6EF9,
32'hBE44A9F2,
32'h3E9284D0,
32'h3E012FBB,
32'hBE8E3691,
32'h3DD81221,
32'hBD6EE0B4,
32'hBE5F7177,
32'hBFBF10F2,
32'h3DA6E19C,
32'hBE890F80,
32'h3E597575,
32'h3E59E355,
32'h3DE163E0,
32'h3E0D0E56,
32'hBEDEEBDB,
32'h3E0EA592,
32'hBC8C9E87,
32'hBE5D6D22,
32'h3DF42224,
32'hBEC86522,
32'hBE475518,
32'h3E9A35BC,
32'hBF2668D6,
32'hBF23AE22,
32'hBF4C93E3,
32'h3CE27019,
32'hBDCF2B40,
32'hBE3C4E60,
32'hBF3F7D5B,
32'h3D246A3F,
32'hBE24AA4B,
32'h3E0E8714,
32'h3EB2D46C,
32'hBEB7E3CF,
32'h3E2E243A,
32'h5DF0FE4D,
32'h3DD09A58,
32'hBF713E44,
32'hBCC9BA35,
32'h3DCF2FBE,
32'hBD5264DC,
32'h3E9063AA,
32'h3E24278E,
32'hBED42AFA,
32'h3E9B57E9,
32'h3EAE2F8B,
32'h3E478F5E,
32'h3E67C4F1,
32'h3CC8D976,
32'hBF8B982B,
32'hBE0A2107,
32'h3E6D19F6,
32'hBEF7C801,
32'hBECC1EF5,
32'hBF413770,
32'hBCC1535D,
32'h3D73DD07,
32'hBF3B6028,
32'hBF3BD941,
32'hBE91AFFD,
32'hBD3AE793,
32'h3DE2C406,
32'h3EAD6007,
32'hBF01DC0A,
32'h3E2CAF34,
32'hBCFCDF26,
32'h3E228004,
32'hBFE94F30,
32'h3D8CC942,
32'hBDDEB21C,
32'hBD42B083,
32'h3E908014,
32'h3E2C080C,
32'hBF739E61,
32'h3DA7C2FA,
32'h3FB12FC6,
32'hBE37174D,
32'h3E3D96E5,
32'h3D01908B,
32'hBFD40A08,
32'h3C7295C4,
32'h3E3F4E8C,
32'hBEBCDE82,
32'hBC71CD47,
32'hBE93A5CF,
32'hBD8CD86D,
32'hBD6C9783,
32'hBF9BC193,
32'hBF3A73BA,
32'hBC9256EC,
32'hBC62CFF0,
32'h3D836BE5,
32'hBEA50E87,
32'hBE8A6A43,
32'h3D9BDF77,
32'hBEC4CEDD,
32'h3D871FB9,
32'hBFB448F8,
32'hBC42783C,
32'hBD6A424E,
32'hBDE908FC,
32'h3DE6C77C,
32'h3C8C64FE,
32'hBEFD456E,
32'hBE8CF416,
32'hBE625D2E,
32'h3E0DEA67,
32'hBDC9ABFF,
32'hBE5FD4A1,
32'hBFCDF6C8,
32'hBF0594F6,
32'h3CA0AD4D,
32'hBF67CE88,
32'h3E1BA67D,
32'h3E019B96,
32'h3CD2C168,
32'hBC7A3E63,
32'hBFFF06DE,
32'hBF341D5F,
32'hBF110111,
32'hBCD5AFE1,
32'h3E4D4570,
32'h3EE251E4,
32'hBE5D9A46,
32'h3E1AE943,
32'hBDAFAF88,
32'hBE30B40D,
32'hBDC7A7D2,
32'h3E3D8EB3,
32'hBE15BBDE,
32'hBECF2C03,
32'h3E1B74D5,
32'hBE983180,
32'hBF14C955,
32'hBDC0AA1C,
32'hBF8E15C5,
32'h3E7C6C68,
32'hBED1B56C,
32'hBED7ABCB,
32'hBFB06B35,
32'hBE6DF559,
32'hBD91B3B8,
32'hBE2D9A81,
32'h3EB4A115,
32'h3E71C463,
32'hBC56D157,
32'h3D2F0476,
32'hBFF2C84E,
32'hBE71EC33,
32'hBD6AD431,
32'hBE9E6828,
32'h3E073358,
32'h3E1243A9,
32'hBE034B94,
32'hBDF0A3CA,
32'hBEC410CA,
32'h3D684DEA,
32'hBFE27E4A,
32'h3DAF9912,
32'h3E87F448,
32'hBECBFD60,
32'h3E914803,
32'hBD8DD2B3,
32'hBEE6B97F,
32'hBF084955,
32'hBFB327D3,
32'hBE8B8EA3,
32'h1755CB82,
32'hBF807B1B,
32'hBFD185C8,
32'hBE727813,
32'hBE9DE172,
32'hBE708926,
32'h3DD6BECA,
32'hBF1958DE,
32'hBD8E5848,
32'h3D2DFF0E,
32'hC00ECFD9,
32'hBEE5D5EA,
32'hBE26ACC0,
32'h071ABA3,
32'h3ED0EF31,
32'h3E9F3322,
32'hBDFF14A6,
32'hBF1EF187,
32'h3CBEA0AB,
32'h3E89C898,
32'hBFA3C723,
32'h3D2F4D3C,
32'hBF2F02C6,
32'hBF4325C3,
32'h3E4B932B,
32'h3E0631D3,
32'hBEB20DED,
32'h3F0CEDBE,
32'hBFAC7641,
32'hBE037FD2,
32'hBE4DCBAE,
32'hBFA640E3,
32'hBF813E5C,
32'hBE00CD8A,
32'hBE3DA659,
32'hBF9B7BBD,
32'hBF44F8AD,
32'hBF17F4DE,
32'h3D70AF93,
32'hBD1670C9,
32'hBFF356D0,
32'hBF1CF13E,
32'h3F05B9D6,
32'h3E289E8E,
32'h3E5EDD36,
32'hBE72597A,
32'hBC857852,
32'hBEE493C5,
32'hBD80EDE5,
32'h3E849EBD,
32'hBF92B233,
32'h1DF21005,
32'hBF18EB18,
32'hBF5FBD18,
32'h3DA81706,
32'h3DCFD55D,
32'hBEC2203C,
32'h3EB11EC9,
32'hBF8532E4,
32'h3E7BCB3F,
32'hBE331D07,
32'hBFBCEABD,
32'hBE6706A9,
32'hBF77C212,
32'hBDA4A43B,
32'hBF60E32F,
32'hBE9BBE69,
32'hBF2B750D,
32'hBC763626,
32'hBC48982E,
32'hC000D23A,
32'hBEBB0EDE,
32'h3E53F2BA,
32'hBC22B865,
32'h3E8F989C,
32'h3DAFBD28,
32'h3E45A151,
32'hBDE21AAA,
32'h3E4AFB0D,
32'h3E04681E,
32'hBF407A7A,
32'hBECA5171,
32'h3E547F56,
32'hBDCD72CE,
32'h3DFED232,
32'h3ED0DE96,
32'hBEF3BB86,
32'h3DBF61FD,
32'hBE85F68D,
32'h1DC08040,
32'h3F71239D,
32'hBFB0BE59,
32'hBDB10320,
32'hBFCBF6E9,
32'h3DE2919F,
32'hBD141497,
32'hBE8A89A8,
32'hBF903FDE,
32'h3D343163,
32'hBC6CEEF6,
32'hC0122DAF,
32'hBE69611C,
32'h3FA19E0F,
32'h3EC7C506,
32'h3F5E6774,
32'h3ED3572E,
32'hBE358657,
32'hBEBE2AB4,
32'h3F78F019,
32'h3EA785C8,
32'hBEC18DD5,
32'hBE238ED0,
32'hBF37BD17,
32'hBFA370C8,
32'hBDBC72A1,
32'h3EC5BEBE,
32'h3DD8743A,
32'hBDBCE314,
32'h3E9F7567,
32'h3D3B8B8E,
32'h3F90C19C,
32'hBF95E9CC,
32'h3E4C443D,
32'hBE80D3EA,
32'h3F2F5718,
32'hBCCE5F04,
32'h3DA978A4,
32'hBF1ACDAF,
32'hBD465BF1,
32'h3CE4342E,
32'hBF11D809,
32'h3E9E0FCA,
32'h3F11840F,
32'hBE1C1BC4,
32'h3F18C495,
32'hBE35C6C9,
32'hBD46543F,
32'hBEA62B83,
32'h3F423E7D,
32'h3F005CCC,
32'hBECBD441,
32'hBE2FBCA3,
32'hBEA99652,
32'h3DE464DE,
32'h3E90690E,
32'h3F342FF2,
32'h3E55B52A,
32'hBF2B83AF,
32'h3F135815,
32'hBFA5D7E3,
32'h3F013379,
32'hBFCD9403,
32'h3EFA98B1,
32'hBF1757B1,
32'hBF1AC88F,
32'hBEE99481,
32'h3DB31272,
32'h3F2005C5,
32'h07587A9F,
32'hBC82FC49,
32'hBF5D0FDF,
32'hBFC9AA40,
32'h3F0DE197,
32'h3E940F64,
32'h3F6847A4,
32'hBE9C8E67,
32'h3F2AD3F9,
32'h3E5FA158,
32'h3EE6EBDC,
32'h3E22E76C,
32'hBEF6FAAB,
32'hBEFB2446,
32'hBCFC83F4,
32'hBEDBEC97,
32'hBD3FEC0B,
32'hBD1AE832,
32'hBEB64174,
32'hBF016B3B,
32'h3EF6B9B4,
32'h3DE99BEC,
32'h3FAED4AA,
32'hBE0E7005,
32'h3F00B54A,
32'hBF08B5B3,
32'h3CB18B03,
32'hBEB4F1BB,
32'h3F403D57,
32'h3ED5B8FA,
32'hBD99A514,
32'h1DCCBA07,
32'hBEB09F07,
32'h3F8B0086,
32'h3FBA0E4A,
32'hBF23E7A0,
32'h400E6E08,
32'hBF8B549D,
32'hBFA39CA5,
32'hBF64C9F4,
32'hBF22386F,
32'h3EB523B3,
32'hBCC41EC8,
32'hBEB6A106,
32'h3FA08A51,
32'h3F21DA02,
32'h3F6F2F5B,
32'hBF17EC9A,
32'hBD0313E1,
32'hBE9B6128,
32'hBD3982DB,
32'h0ED962E8,
32'h3F7E01B2,
32'hBE1F9869,
32'h3F602471,
32'h3E8C2E48,
32'h3E1A43EA,
32'hBD9DB51D,
32'h3EAF1BA4,
32'h3E966D91,
32'h3C81BC53,
32'h3DAB5963,
32'hBF1BF8E1,
32'h3F5AC266,
32'h3F22A7BF,
32'h3E8F0000,
32'h3C2BF94B,
32'h3E2DD71A,
32'hBE7578F0,
32'hBDDC217B,
32'h3F7C180B,
32'hBF34FB2E,
32'h3C9FF29B,
32'hBF1861D9,
32'h3F5C0ECF,
32'h3F0A3E14,
32'hBE82CA4B,
32'h3D4BAE31,
32'h3D0BC5D7,
32'h3D89CBAA,
32'hBDD95C02,
32'h3DB8E889,
32'h3F3DD4BA,
32'h5DF45D00,
32'hBD96314C,
32'h3E41CE16,
32'h3D254D01,
32'hBC0772D1,
32'h3D032D97,
32'h3E9B952B,
32'hBCA714FF,
32'h3D372778,
32'hBCDAA203,
32'h3F5819E6,
32'h3EF044FE,
32'h3E8CAF16,
32'h3D95442A,
32'h5DF53C97,
32'hBE95BC30,
32'hBCBE3148,
32'hBDF1463C,
32'hBF01490E,
32'hBCC627EF,
32'hBF698331,
32'h3F639A63,
32'h3CD90497,
32'h3F215CC3,
32'hBE84C375,
32'h0EDD4C14,
32'hBD35CA4A,
32'h3DDF30B3,
32'hBD945680,
32'hBD20C924,
32'hBC10EFF6,
32'h3D5CB4A1,
32'hBCFF58D8,
32'h40800013,
32'h2ED40212,
32'h3CBEF4D1,
32'hBD8545DF,
32'h3CE2B0D9,
32'hBC1FD474,
32'hBD62DAFD,
32'hBDA044CA,
32'hBD34A3B7,
32'h3C3EC657,
32'hBCE87816,
32'h3C9A34C4,
32'h0EC78535,
32'h1DF01AE3,
32'h3DB5D201,
32'h3D66911A,
32'h3C868D44,
32'h3D81F071,
32'h5DF54391,
32'h0EC45377,
32'hBC6CC889,
32'h3D6D4964,
32'h5DEEB417,
32'h3D919C82,
32'h3CA362D0,
32'h1DD55CCB,
32'hBC7DDF6D,
32'h3D1FA427,
32'h3C80CFF7,
32'h3D2DD121,
32'h3CCD4FE7,
32'h3C755C32,
32'hBC5158A4,
32'h3C0EFD12,
32'h3CCDD566,
32'hBCC9DBB5,
32'hBD6CE35C,
32'h3D9D5CC3,
32'h1DEB8B43,
32'hBCA67C58,
32'hBD6FD832,
32'h3C73600E,
32'h3D247BFE,
32'hBCEE8503,
32'hBDC03513,
32'h5DF5D49E,
32'hBCF7A08D,
32'h3D392CC3,
32'hBD83036D,
32'h5DC8B2A0,
32'h3D0DAAA1,
32'hBD38F52D,
32'h3DAC646F,
32'hBCB069E2,
32'h3D2DEC07,
32'h3C91AA34,
32'h0EC391F3,
32'hBC2A2151,
32'h2EDFAA66,
32'h3CF16379,
32'h3D19AFE1,
32'h5DF4F81D,
32'hBC4C2564,
32'hBC385DF8,
32'hBA092CE,
32'hBD8731DA,
32'h3D8F95CB,
32'h3D78090C,
32'h3CC1470F,
32'h3D928D01,
32'hBD4D35BD,
32'h3D8026B9,
32'hBD00281A,
32'hBCF8551F,
32'hBC31625F,
32'h3D3CF997,
32'h3DAE89E7,
32'h3DC54422,
32'h3DA941B3,
32'h3D0A1420,
32'hBCB0BB93,
32'hBD99154A,
32'hBCC4D46C,
32'h1DD50A44,
32'hBCDC78E7,
32'h3E1B0194,
32'hBD56DD01,
32'hBD6EE40E,
32'hBCF41605,
32'hBE12E45A,
32'h3EA63A68,
32'hBD12184A,
32'hBCAB3023,
32'h3D64E10D,
32'h3CC50F96,
32'h3CAD5FF3,
32'hBD996C16,
32'h3DD8E604,
32'hBDD8E1F8,
32'h1DEC7620,
32'hBDA6019B,
32'h3D48DEC1,
32'h3F13EEFF,
32'hBEBAD3DA,
32'h1DC35538,
32'h3E171A82,
32'h3CEA3088,
32'hBF4F833E,
32'h3E95132D,
32'hBDDE5F9C,
32'h3EC8FF7C,
32'h3D64B347,
32'hBCA900CE,
32'hBCAADB2C,
32'h3DFA9C7E,
32'hBC80DD36,
32'h3DF43D07,
32'h3D500DE7,
32'h3F937DB1,
32'h3EBFAC85,
32'h3C031ABD,
32'hBE9F9860,
32'hBE2FF308,
32'hBCB49DC3,
32'hBC9813E0,
32'h5DFE4E20,
32'h3C15CEAB,
32'hBDDBA05F,
32'h3CA96F62,
32'hBE9FD89B,
32'hBE49952B,
32'hBCB395BF,
32'h3E645DFF,
32'h3D47D123,
32'hBD0F6770,
32'hBED87F39,
32'h3DD7AE0F,
32'hBD7FA677,
32'hBDDBD0B5,
32'h3F426F5B,
32'hBF314BC6,
32'h3E03F3FB,
32'hBD1C6A9F,
32'hBE0BB568,
32'hBF194A7C,
32'h3F6FA6DF,
32'hBEE625EF,
32'hBE9F01C9,
32'h3F7154D8,
32'h3D81518A,
32'h3FDB690E,
32'hBE988BDE,
32'hBD49C528,
32'h3C45B1EE,
32'h5CC2D54,
32'h075988C0,
32'hBE53E12E,
32'hBE50C3F4,
32'hBEC9484D,
32'h3F1CE9FD,
32'hBF5E421C,
32'hBED2DB9D,
32'hBEF1093A,
32'h0ECDBE30,
32'hBF366225,
32'h3EEF88C7,
32'h3D145E26,
32'h3E218430,
32'h3F0297F8,
32'hBDA4D108,
32'hBEA45ECE,
32'hBE123FDC,
32'hBDE78868,
32'h3E266D27,
32'hBE81D765,
32'h3E9247AD,
32'hBF7F9539,
32'hBDEC9D77,
32'h3F3EEB06,
32'hBE564BD7,
32'h3F3E75F2,
32'hBE5332B5,
32'hBE231709,
32'hBE0DDD69,
32'h3DBD0CDA,
32'hBDB0D4FB,
32'hBFAC18AB,
32'hBF941ADC,
32'hBE5B7F63,
32'hBE6A54BD,
32'hBF9DB401,
32'hBF3E87EC,
32'hBE96D47B,
32'h3D8CDF3A,
32'hBF7222BA,
32'h3F096E30,
32'hBC933A4A,
32'h3F14377D,
32'h3E575548,
32'hBF7AFC14,
32'h3E0210CE,
32'hBE122875,
32'hBE829BAB,
32'h3E09FF04,
32'hBE97BE1F,
32'h3EB8AA18,
32'hBE434060,
32'hBED8AFAA,
32'h3E02A9F7,
32'hBE953588,
32'h3EDBA8BB,
32'h3D12A838,
32'hBF4241D9,
32'hBE404233,
32'h3D6FDED4,
32'hBD20EF0F,
32'hBFC1DDE9,
32'hBF5F61C1,
32'h3EFEFD0A,
32'hBF02DE67,
32'hBFACDABB,
32'hBF0A98F7,
32'hBF482D65,
32'h3E707772,
32'hBF43B326,
32'h3F0B6199,
32'hBD0971DB,
32'h3F72C8B9,
32'h3ED56688,
32'hBEAC201A,
32'h3F2ACE67,
32'h3D8953F4,
32'hBE992881,
32'h3DCC7547,
32'hBCE8C162,
32'h3E85FBAE,
32'hBCAE01CA,
32'hBE658193,
32'h3EECA8F0,
32'hBF24B3E4,
32'h3F20981F,
32'h3E6F1BE1,
32'hBF13389C,
32'hBEAC5CBE,
32'hBD1921F4,
32'hBD8A40B8,
32'hBEE6C305,
32'hBF6A9A27,
32'h3F427BDD,
32'hBEDF0C8E,
32'hBF8285D0,
32'hBF1473D4,
32'hBEB71937,
32'h3F361425,
32'hBF104655,
32'h3F6C3897,
32'h3C04A5A8,
32'h3F1D2722,
32'h3E981452,
32'h3E4A8056,
32'h3F1F64D1,
32'hBCEAAE4A,
32'hBEE4E20D,
32'hBF6181C2,
32'h3F03244C,
32'h3E0958DF,
32'h3EEA0393,
32'hBF54A40B,
32'h3F0C9682,
32'hBEAA3273,
32'h3F4109DF,
32'hBF5A3F19,
32'hBF098D84,
32'hBDE8035C,
32'hBD97D008,
32'hBC01CC32,
32'hBCAE9512,
32'hBFAC54B7,
32'h3F1AF9EA,
32'h3DAD23B0,
32'hBE71ECBE,
32'hBED0D7AE,
32'hBD96D6DF,
32'h3E2D58DD,
32'hBEC98225,
32'h3F0746B0,
32'hBCBCC13D,
32'h3D7B1188,
32'h3EF80343,
32'h3EAC3036,
32'h3EF4AC76,
32'hBEBD3B40,
32'hBF35F8E6,
32'hBF39152E,
32'h3E5C7CF0,
32'h3E92045A,
32'h3E025C43,
32'hBF83FD70,
32'h3D51081B,
32'h3DE9C089,
32'hBEB4D92E,
32'hBFD99396,
32'hBFC05053,
32'hBE0ABAA3,
32'h3D7D5AC8,
32'hBC7144AC,
32'hBFE79AF7,
32'hBFAEC2AB,
32'hBEB558C0,
32'hBE22C984,
32'hBE0ED296,
32'hBECF0456,
32'h3DB40FCB,
32'hBF93781E,
32'hBDBD25BB,
32'h3F3223EF,
32'hBD1AB9D0,
32'h3E60F4AF,
32'h3E111CFA,
32'h3E7BAB1C,
32'h3EF5E529,
32'hBDE63C59,
32'hBF192A8C,
32'hBF787246,
32'hBCB65291,
32'h3E82D3CE,
32'hBD076222,
32'hBF9AAD12,
32'h3D6ADF9A,
32'h3E3363D7,
32'h3EFD9F22,
32'hBF0E59B5,
32'hBF789515,
32'hC00DA2BA,
32'h3D8F2A91,
32'h3CC25AEE,
32'hBF84453B,
32'hBFA2A1F6,
32'hBF7773EC,
32'hBE4082C2,
32'hBF774A9A,
32'hBE7132D6,
32'hBEC7541B,
32'hBEACFDC1,
32'hBE2B33E2,
32'h3EF2DB30,
32'h1DFFCDE6,
32'h3EC47DA8,
32'h3E6DCD38,
32'hBE0CEB92,
32'h3EC06A3C,
32'h3E7EE1EA,
32'hBE988B40,
32'hBF523800,
32'h3E9413BB,
32'h3E9AF6A1,
32'h3DE00CD8,
32'hBFAFAE37,
32'h3ECE8386,
32'h3DD2C839,
32'h3DCB1553,
32'h3DAAA721,
32'h3EBCAA5C,
32'hBFF6DA39,
32'h3D8B6FF5,
32'h3D10251F,
32'hBFB27586,
32'hBF7DD6C3,
32'hBEFF0E09,
32'hBEAA3B6F,
32'hBF7CB63A,
32'h3D235B76,
32'hBE38ABFF,
32'hBEA918B2,
32'hBEC09CCF,
32'h3E8ADC07,
32'h3E803700,
32'h3E20BB5A,
32'hBD4C3622,
32'h3CC77128,
32'h3EA04ED3,
32'h3C97625A,
32'h3D0601C8,
32'hBF41FAF4,
32'h3E3E58A3,
32'h3E7B69F0,
32'h3EE92EC2,
32'hBF62CFE6,
32'h3E0A8C42,
32'h3F1E6ABC,
32'hBE729F17,
32'h3D7CB945,
32'h3E8B37C1,
32'hBFE8D801,
32'hBDB1A30D,
32'h3C8444FC,
32'hC0072126,
32'hBF5AED2B,
32'h3EE6CB93,
32'hBEB66E0E,
32'hBFA85B55,
32'hBCE05124,
32'hBCA888AD,
32'hBE934493,
32'hBE8EB051,
32'h3E1B93B8,
32'hBE2BCD10,
32'hBE9EC7ED,
32'h3E4E0DF7,
32'h3E98633A,
32'h3E9BB89A,
32'h0ECB4538,
32'hBED47EB1,
32'hBFC80221,
32'h3DC48BC8,
32'h3C40721D,
32'hBDB13535,
32'hBFAC862B,
32'hBF56ACCE,
32'hBEB4B002,
32'h3F066309,
32'hBE1C5307,
32'hBE8CD2A1,
32'hBF5E0147,
32'h3D7EE954,
32'h3CCA560B,
32'hC0010B8B,
32'hBF72BF3C,
32'h3EAE72A1,
32'hBD01C4C4,
32'hBEE45BCC,
32'hBED8209F,
32'h3D2C715B,
32'hBE634B4D,
32'hBD9829E5,
32'h3E8CA50E,
32'hBF097B5F,
32'hBE8E43C8,
32'hBE26531A,
32'h3D6DA1FC,
32'h3EDE6B97,
32'h3D95CF15,
32'hBF1DE47C,
32'hBEFF63D7,
32'h3EB32D75,
32'h3ECAE50D,
32'h3E65A70C,
32'hBFC21999,
32'hBFD6FD8E,
32'hBEA037E9,
32'h3E9186DE,
32'h3E8BEE6F,
32'h3C5B428E,
32'h3E9013A4,
32'h3D8B5B12,
32'hBD75E76C,
32'hBFEB588B,
32'hBF84E5C8,
32'h3E667657,
32'h3D047B5B,
32'h3E18EB85,
32'hBE137073,
32'h3DD3CA7F,
32'hBEB4A187,
32'hBD4F7330,
32'hBC0A9241,
32'hBF337791,
32'hBE1853F6,
32'hBEC85CC8,
32'h3DF61D09,
32'h3E439FEB,
32'h3D929A56,
32'hBE90C38C,
32'hBF53BEAA,
32'h3C2A585A,
32'hBE1A776A,
32'h3ED58944,
32'hBF75E037,
32'hBFF9F36D,
32'hBDE82108,
32'hBEA92C89,
32'h3EAA0E80,
32'hBDB27081,
32'hBF72602A,
32'h3D558510,
32'h3CAED09B,
32'hBFC67C46,
32'hBFFE0AB9,
32'hBF398235,
32'hBE9E690D,
32'h3F369B91,
32'hBE00A4F7,
32'hBD434C91,
32'h3E7D66C5,
32'h3C9CA322,
32'h3E5F26F3,
32'hBE88D5C6,
32'h3EF65DA6,
32'hBEA0DB5B,
32'h3E97D67D,
32'h3EDC5CC3,
32'hBD546E6B,
32'h3EB4F68D,
32'hBF31D4FD,
32'hBF6A1D8E,
32'h3E9D18E9,
32'h3E846445,
32'hC023E397,
32'hBFD043E0,
32'hBF07DDC8,
32'h3E87368A,
32'h3CD12743,
32'h3E94594E,
32'hBFDB0055,
32'hBCFEC3F2,
32'hBDA75260,
32'hBFA07711,
32'hBF67B591,
32'h3E3017BC,
32'hBE2DF59B,
32'hBF0821B6,
32'hBEE3021D,
32'h1DDE5E63,
32'hBE8C037A,
32'hBEF69534,
32'h3EA777A2,
32'hBF517278,
32'h3E99057C,
32'hBE1D23EB,
32'h3EE066BA,
32'h3ECA0410,
32'hBE8056FE,
32'h3E7A5AED,
32'hBF9EFAC5,
32'hBF1D9039,
32'h3E8B42CF,
32'hBE2EF522,
32'hC030D317,
32'hBED4AA3E,
32'hBEB941EB,
32'h3E570C42,
32'h3DD292CC,
32'h3E14721B,
32'hBF83B623,
32'hBA0B660,
32'hBD2BEE81,
32'hC01371BA,
32'hBEBF2F21,
32'hBE9FA3FF,
32'hBA50135,
32'hBF1C3F89,
32'h3E8B2D00,
32'hBE5C6CA5,
32'hBEA4B6F4,
32'hBEBE8AEE,
32'h3F63675A,
32'hBDECBE49,
32'h3D884519,
32'hBE8F5DCB,
32'h1DDE5F5D,
32'h3E8DF759,
32'h3F3D5684,
32'h3F127284,
32'hBF7EB247,
32'hBF356C91,
32'hBE8ACA12,
32'hBEE10498,
32'hC0299AD2,
32'h3E192119,
32'hBF6AC04A,
32'h3EB2BA6D,
32'h3E6A3A3D,
32'hBED1979A,
32'hBF44E646,
32'h0EC64634,
32'h3D8FFEB0,
32'hBFFDF40F,
32'h3EC35913,
32'hBE6755CF,
32'h3EA2E0C4,
32'hBF016787,
32'h3E650E70,
32'h3E50F770,
32'hBF303A1A,
32'hBD6E0DC3,
32'h3E95C0E5,
32'hBD07E8C7,
32'hBDF9183D,
32'h3DC906CF,
32'h3E971BDD,
32'h3E016FC1,
32'h3F1F445B,
32'h3F0E2D82,
32'hBEE29437,
32'hBEEC7848,
32'h3F2295AA,
32'hBE88ACA6,
32'hC02D1877,
32'hBEC0AA46,
32'hBF3AD8E5,
32'h4008CE63,
32'h3EF6EFAC,
32'hBE52C25D,
32'hBEE656C0,
32'h3C97A888,
32'hBC0E60EA,
32'hBFEFA501,
32'hBEC0945C,
32'hBE67214D,
32'hBECF42A5,
32'hBEEF0144,
32'hBEDC1CA7,
32'hBE9D18B4,
32'hBEC7A153,
32'hBF0AB76C,
32'h3E6F9DF9,
32'hBF55BF3B,
32'h3EB62415,
32'h3E835FFF,
32'hBEA8A5A0,
32'h3F437FD9,
32'h3EBD9B95,
32'hBE01DCAB,
32'hBFD544D5,
32'hBE1C7546,
32'h3EBA4DF6,
32'hBE9B502E,
32'hBFB886BB,
32'h3EB80A00,
32'h3E4256EE,
32'h3E1A08DB,
32'h3F374716,
32'hBE17B5D9,
32'hBED65C5E,
32'hBCA50CD2,
32'h5DC4DCF4,
32'hBF9FF2B5,
32'hBF84C6F0,
32'h3ED3972A,
32'hBE09D4E5,
32'h3F48B3E2,
32'hBEED0E39,
32'h3C293177,
32'hBF20737D,
32'h3EDF976C,
32'hBE081091,
32'hBDF7CCA9,
32'h3EB6F073,
32'h3EA57CE3,
32'hBF85EE23,
32'h3D1FE944,
32'hBE524D07,
32'hBE7834EA,
32'hBFB602C7,
32'hBE41108E,
32'h3F404741,
32'hBEE658AD,
32'hBF658380,
32'hBE499945,
32'hBDD4B401,
32'hBEDB8BE4,
32'h3F213077,
32'hBEBC6F9D,
32'h3D9D08EB,
32'hBCF2C644,
32'hBDB59A44,
32'hBFC0E6DE,
32'hBF84221F,
32'hBD6AF31D,
32'hBF084E77,
32'hBE86D2A7,
32'hBF243D79,
32'hBEA2BB7B,
32'hBEF59084,
32'h3DF1216C,
32'h3EE14FED,
32'hBCD10B5C,
32'h3F06885A,
32'hBF0FFC14,
32'hBF947612,
32'h3D1BA11C,
32'h3E98556E,
32'hBEE100AF,
32'hBFCC6D22,
32'h3ECF0D1D,
32'h3DABC70F,
32'hBFA0F7B1,
32'hBF7B6849,
32'h3D5B8C48,
32'hBE2138BF,
32'hBF1FEC49,
32'h3F22FA23,
32'hBEE9BA15,
32'h3E273399,
32'hBD0EB3FA,
32'h0750C39E,
32'hBF562165,
32'hBF268D17,
32'hBD9FCF40,
32'hBF8ABD27,
32'hBE1A014D,
32'hBE6BDEBF,
32'hBF8A019D,
32'hBF819FA5,
32'h3EC05931,
32'h3F7E2BF2,
32'hBD642556,
32'h3F3902C6,
32'hBF6D06E2,
32'hBF30B481,
32'h3E2BF09C,
32'h3EF1B30F,
32'hBE5BC09A,
32'hBEFCDA1C,
32'hBF988F12,
32'hBEBDCBA3,
32'hBF8B247F,
32'hBF9DE506,
32'h3CEB0280,
32'hBF0B43AA,
32'hBF87F607,
32'hBF91A9A1,
32'hBE71DF6C,
32'hBD807E7B,
32'hBD3DE63B,
32'h0EDCF531,
32'h3F014463,
32'hBE053EB8,
32'h3E71D77D,
32'hBF8B9A74,
32'hBE463C69,
32'h3ECA94F8,
32'hBE2AC428,
32'hBE8EE758,
32'h3F8F663A,
32'h3F149B96,
32'hBD647DD6,
32'h3DB5ACB5,
32'h3E94FC02,
32'hBEA8AAF2,
32'hBF815633,
32'hBD972DA8,
32'hBD9FB4F4,
32'h3E4E5825,
32'hBDB38B16,
32'h3D3031AA,
32'hBF095380,
32'hBEC0F227,
32'hBEBB5730,
32'hBCD46E81,
32'hBC33FE8F,
32'h3D07E7CE,
32'h3D7A9904,
32'hBDDBCDAC,
32'hBD279A48,
32'hBD34CBCD,
32'h3E12A0A7,
32'h3F3B8699,
32'h3F052693,
32'hBFC69B81,
32'hBC6542D3,
32'hBE8DDF78,
32'hBEF1C108,
32'hBF3B89E0,
32'hBE9AB116,
32'h3FBCA836,
32'h3C826799,
32'hBE3D3BE4,
32'h3ED01D5E,
32'h3EE4E7A7,
32'h3EAF1204,
32'hBE2056D1,
32'hBD7AF515,
32'hBF3A6748,
32'hBD154714,
32'hBC944C02,
32'h3E9ED049,
32'hBD9CA709,
32'h2EDF8415,
32'hBD618C43,
32'hBDB0D2A7,
32'h3D53E21D,
32'h3DC0D87D,
32'hBD32AB10,
32'hBD22563E,
32'hBD87A0F1,
32'hBD5931A9,
32'h3F485634,
32'h3EF41EE1,
32'h3E324D19,
32'hBC893770,
32'hBDC377AA,
32'h3F098106,
32'hBDC5A2B9,
32'hBD99699A,
32'hBF5CAF5C,
32'hBCB986BB,
32'hBEA01876,
32'h3F0BC358,
32'hBDB8EE6E,
32'hBE32D889,
32'hBD6FD9DD,
32'h075B5BEE,
32'hBD9015F2,
32'h3D2A1BAA,
32'h3DE40D70,
32'h3F3D923D,
32'h3D8C6A3D,
32'h3CE56783,
32'h1CEE014,
32'h3D9E859B,
32'hBC870B8B,
32'h3DA18B79,
32'hBD505769,
32'h3D0C4387,
32'h3D7F0C1C,
32'h3D2D53E0,
32'h3F5C7456,
32'h3F1CC153,
32'h3E85C4CB,
32'h3D83555F,
32'h3C944F0C,
32'hBEAF7C88,
32'h1DC191D4,
32'hBD7A75BB,
32'hBE89D04B,
32'h3C51AA99,
32'hBF50C76D,
32'h3F42C41C,
32'h3D8AC586,
32'h3F2F5718,
32'h3D5F865E,
32'hBD73A8E3,
32'hBDB8966B,
32'hBD81AE7A,
32'hBD888D49,
32'h3DBFDBBC,
32'h3D266DB0,
32'hBCA0FE22,
32'h17548C55,
32'hBD2D87B6,
32'hBC06C34A,
32'h3D8F684E,
32'hBCD8CCA3,
32'hBA6DB97,
32'hBD13F4EA,
32'h1DDBA822,
32'h3DB74AF5,
32'hBD3F3854,
32'h5DF407EB,
32'h3D33D8E6,
32'h3D74DA87,
32'hBD460F5C,
32'hBCB7D226,
32'h2EC6617C,
32'h3D3C54BC,
32'hBD98F8B0,
32'h5DF00B02,
32'h3CA6A36D,
32'hBD6501FD,
32'hBDE16B65,
32'h3CBEA477,
32'h1DC40FFF,
32'hBD6F0AC0,
32'hBDA1A6F9,
32'h3D6767E2,
32'h3D9AC9DA,
32'hBC1AF644,
32'hBDAF2D57,
32'hBDAB6435,
32'h3D788EAB,
32'h3DB610FF,
32'hBDA337A1,
32'h3D3B6AE3,
32'hBD4702EC,
32'h3C247AA8,
32'hBD2212C0,
32'h3D4757F5,
32'h3D7DBC1D,
32'h3DD544EE,
32'hBC2D6593,
32'hBDC43455,
32'h3DDC9DD6,
32'hBD46CA92,
32'hBC84A6A9,
32'h3D89DDF2,
32'hBD22A905,
32'hBCAB70EA,
32'hBC05E09F,
32'hBC85D592,
32'hBD36BD71,
32'h3D82D3BA,
32'h3D1B7975,
32'h0EC2D62B,
32'h3C8F1C36,
32'h3C6DD145,
32'hBD738837,
32'h0755698B,
32'h3D754B2B,
32'h3CB9AE98,
32'h3D0D537E,
32'hBC825B7F,
32'hBD18D327,
32'h3DA626D3,
32'hBC900068,
32'h3D0BB5E6,
32'h3C63AB51,
32'hBC8ED068,
32'h3CBEF4A5,
32'h3DBAE513,
32'h075BED0F,
32'hBC55DFFD,
32'hBC933608,
32'h3D901562,
32'hBC7013DD,
32'h3D35EC40,
32'hBD81AA01,
32'h3D8D00BC,
32'hBD7A5F91,
32'h3D9B5407,
32'hBC5AC818,
32'h3D76EBAC,
32'hBD0C95AC,
32'hBD4351B2,
32'h3D302D95,
32'h3D8F1D3E,
32'hBCC7035E,
32'hBCB1322C,
32'hBD0369BF,
32'hBCFE3715,
32'h3DE4EEC8,
32'h3CE71E8F,
32'h2EDA0965,
32'hBD56355B,
32'h3CE7186E,
32'hBC73EC8D,
32'h3D219F17,
32'h1DC86AE4,
32'hBC4465F3,
32'h3D201D51,
32'h3D7CED06,
32'hBC5F1592,
32'hBD34666C,
32'h3D31CEB8,
32'h3D3BB199,
32'hBDB0F264,
32'hBD203717,
32'hBCC8C3D1,
32'h3D6912D7,
32'h3D2B07D2,
32'hBD791259,
32'h3CC423FF,
32'hBD8CDE58,
32'hBCBFD288,
32'h3D90A916,
32'h3D3B3999,
32'h3DB12B8E,
32'h3D1A1867,
32'hBC0F6E0F,
32'h3D2E2863,
32'h3C42AAA0,
32'h3C8942DD,
32'h3C48C3F2,
32'hBD994B2B,
32'h3CB1B956,
32'hBD3E0E6F,
32'h3CA62399,
32'h0EDE3A9B,
32'hBD6E6A1E,
32'hBD076574,
32'hBD439329,
32'hBC46D282,
32'h3CBF05DA,
32'h3C230CE3,
32'h3DA3F4C0,
32'h3D63784C,
32'h3DCBF437,
32'hBC751CA4,
32'h5DF69999,
32'h3DB8B5F8,
32'hBD0C1DFE,
32'hBD3CC708,
32'h3CA5343E,
32'hBD9DC4BA,
32'hBD13C7C3,
32'h3F2A8C56,
32'hBF449159,
32'h3CDEBE61,
32'h3EE8970B,
32'hBEABD3E7,
32'hBF1CFEF5,
32'hBF2402A6,
32'h41000002,
32'hBDDC80D0,
32'h3D08FDC1,
32'hBD7920CA,
32'hBDA1D73B,
32'hBD8FE423,
32'h3E5ED5EF,
32'h3F082EE4,
32'hBE403D88,
32'hBEB96455,
32'h3E0B3F2E,
32'h3E238FDC,
32'h3DC91A7D,
32'hBF190442,
32'h3D0FDC9D,
32'h3F2C3447,
32'hBED52706,
32'hBEF404E2,
32'hBE8704DD,
32'h3D2F03F6,
32'hBDBAFC97,
32'h3E97B39E,
32'hBE32153A,
32'hBEA1EEAF,
32'hBF0F6E03,
32'hBEA251FC,
32'h3EDC8C06,
32'hBF31CA56,
32'hBF04E74E,
32'h3E938DB1,
32'h3C9556E0,
32'h3C19D987,
32'h3CD441FA,
32'hBDB68F2D,
32'hBEC0894D,
32'hBDF4A5B3,
32'h3EEDB915,
32'h3DB1576C,
32'hBEBC2001,
32'hBF07EF1D,
32'hBF4E0F00,
32'h3DF94E51,
32'hBEFE057D,
32'hBF003D98,
32'hBD350C0E,
32'h3F6C1C58,
32'h3D672026,
32'hBFAB3C1E,
32'hBF03342B,
32'hBE6798E3,
32'hBE2E4F8E,
32'h3E583EFE,
32'hBECCBCC2,
32'hBE608BD7,
32'hBEC99621,
32'hBEA6F35A,
32'h3ECBFF62,
32'hBE24D063,
32'hBEAC9C4D,
32'h3F3B292C,
32'hBECDDB07,
32'h3E432171,
32'hBD006C06,
32'hBD020FF9,
32'hBF1C1B01,
32'hBC837799,
32'h3EA8C24F,
32'hBE646A0B,
32'hBE022D4F,
32'h3D48CF45,
32'hBEDD448B,
32'h3E5724E7,
32'hBF0C1865,
32'hBE88C2D5,
32'h3D671F5A,
32'h3E5250F2,
32'hBD8DFD36,
32'hBF3CE0C2,
32'hBED05288,
32'hBEB56895,
32'hBD85FE2D,
32'h3E053C65,
32'hBF57A588,
32'h3E235CA9,
32'hBD320539,
32'hBE52DE85,
32'h3F3EA8E4,
32'h3F3B2353,
32'hBF81667C,
32'h3F6D0ADE,
32'h3EA3A43D,
32'h3E5824BF,
32'h3C6BEC75,
32'h3C3220A4,
32'hBFF294BE,
32'h3D943277,
32'h3EB0E041,
32'hBDECF87C,
32'hBEC729A0,
32'h3E5C7B35,
32'h3EB15696,
32'hBC4BA3A2,
32'hBFAC418B,
32'h3EC70B71,
32'h3C26C1F1,
32'hBE9A8A28,
32'h3C7C1EB4,
32'h3F3E5F17,
32'h3EAE4BF3,
32'hBE66E486,
32'h3D38EC1F,
32'hBEC55C9C,
32'hBF8014F2,
32'h3EA25666,
32'h3E0CD120,
32'hBEFABDC4,
32'hBD969CCF,
32'hBEBE2810,
32'h3C91CB7A,
32'h3ED591D8,
32'h3E505ADD,
32'h3E9BFC8A,
32'hBD086D24,
32'hBDA573A6,
32'hBFA5BEDB,
32'hBE3B7634,
32'h3F479271,
32'h3E280288,
32'hBF830505,
32'h3F6F31FB,
32'h3ED2B6F3,
32'hBEF9A8A4,
32'hBF3E8376,
32'h3EA9F3B8,
32'h3C4C8B9F,
32'h3E363A7D,
32'h3EE4785E,
32'h3F335E83,
32'h3E831944,
32'hBF5A7C7C,
32'hBE87B1AE,
32'hBF6ECE4E,
32'hBED4AADF,
32'h3ECDAB49,
32'h3EA8B367,
32'hBFA7CCEA,
32'hBEAAF1FC,
32'hBF01DF5C,
32'h3E24799F,
32'hBE95AC75,
32'hBF6BE9FF,
32'hBDFD2B33,
32'h3D388CB1,
32'h3CA2ABE1,
32'hBF11BCC9,
32'hBF0AA7F0,
32'h3EE3653E,
32'h3E84C5A4,
32'hBF3BE395,
32'h3D04858B,
32'h3FA8FDD2,
32'hBF8DA8BB,
32'hBF78CBC6,
32'h3F01C8CA,
32'h3DC50C26,
32'h3F096B53,
32'hBE7B6871,
32'hBE18E95F,
32'h3E1491A7,
32'hBE91F2A0,
32'hBEED87E3,
32'hBFDCAD34,
32'hBE867152,
32'h3C103F1A,
32'h3F15033C,
32'hBFA1D73B,
32'h3F26F0A5,
32'h3F01D2A4,
32'hBD70460A,
32'hBE4AEBF4,
32'hBF4BB764,
32'h3D72F673,
32'h3C20F1C9,
32'h3D80A903,
32'hBF06FA51,
32'hBEBAA648,
32'h3EB68D00,
32'h3E11D986,
32'hBE3E9345,
32'hBE94C5F7,
32'h3EF80665,
32'hBE91EDDD,
32'hBF3AF38F,
32'h3F1E5E38,
32'h3E9E9C6E,
32'h3ECE046B,
32'h3EACD935,
32'hBF55F830,
32'h3E13C36F,
32'hBEB6DA8A,
32'hBD8F0067,
32'hBFC58E42,
32'hBEA34BA9,
32'h3DB6E257,
32'h3C34924F,
32'hBEFA0317,
32'h3F84909F,
32'h3EDF17D0,
32'hBE49198C,
32'h3F107BF9,
32'h3E326547,
32'hBF010BBF,
32'h1DF9FB64,
32'hBDA2727F,
32'hBF0D2BD2,
32'hBF0A6976,
32'hBF3AFC7C,
32'hBDB71F09,
32'hBF3A9E2B,
32'hBF818E50,
32'h1DCE58C4,
32'hBE11EA07,
32'hBF0A4C59,
32'h3F0B3DB6,
32'h3E10367D,
32'h3F1BAF54,
32'h3EE03F91,
32'hBF4AF6D6,
32'h3F25F653,
32'hBE98EB46,
32'hBE97EF3A,
32'hBF689DEE,
32'hBF576294,
32'hBE09D033,
32'hBE8DD3E1,
32'hBF0D8254,
32'h3E50B7C1,
32'hBF24AD97,
32'h3E30DF2D,
32'h3F40595D,
32'h3E2B8F5E,
32'hBFA5AC49,
32'hBD83E018,
32'hBD96510B,
32'hBEFEBE68,
32'hBE75097E,
32'hBEA178AF,
32'hBE4904F5,
32'hBF32F752,
32'hBEE2EE7C,
32'h3EA49568,
32'h3D76E9B4,
32'hBF66CC68,
32'h3F24D50E,
32'h3E18FA81,
32'h3EF7EE07,
32'hBE07C9C4,
32'hBF19464E,
32'h3EC67CF1,
32'h3D40A9A4,
32'hBDBFD10A,
32'hC01BDA1D,
32'h3F38F976,
32'h3EB82BD1,
32'h3F5CBB69,
32'hBFB74021,
32'h3EF90EB7,
32'h3EE863A7,
32'h3F08E2E5,
32'h3F146855,
32'hBDAA0A60,
32'hBF343495,
32'hBD1BD376,
32'h1CDDA07,
32'hBFA9A76A,
32'hBDEBC7B1,
32'hBEAC471A,
32'hBE66C06C,
32'hBDE9AB65,
32'hBF04B704,
32'h3ECB5E52,
32'hBE26D91E,
32'hBF6DA993,
32'h3F143976,
32'h3DCF59A7,
32'h3F14C286,
32'hBD83E8B6,
32'h3EB0693C,
32'h3F1F14AF,
32'h3F2818F8,
32'h3F120B68,
32'hBF169C4F,
32'hBC8B4360,
32'h3E844F51,
32'h3F1D1F5A,
32'hBF815A76,
32'h3EB2B05F,
32'hBEC6F8CD,
32'hBF713156,
32'h3DAAF335,
32'hBEFD3A32,
32'hBF9DA423,
32'hBD7FF47A,
32'h3D4838E6,
32'hBF98B9E8,
32'hBECB61B4,
32'h3E9CFFD0,
32'h3ED563E5,
32'hBECBB412,
32'hBF284525,
32'h3F10C2C5,
32'hBF593C7F,
32'hBF7BD689,
32'h3E8FC031,
32'hBDA23CE2,
32'h3EF70C80,
32'h3EDF91B1,
32'h3C784EB0,
32'h3E90B34C,
32'hBEBB5DF2,
32'h3E38B7C1,
32'hBF25D5E1,
32'hBEEA2540,
32'h3E9D483A,
32'h3E9389C4,
32'hBF837D01,
32'h3EC7B6A8,
32'hBDB7DBED,
32'hBF9AF458,
32'hBD57CC27,
32'hBF9F6E46,
32'hBF338108,
32'h0ED53DFD,
32'hBD8719BD,
32'hBE714A77,
32'hBEF0EC94,
32'hBE41C542,
32'h3C3F3F60,
32'hBDA75398,
32'hBFAB0C5D,
32'h3D7F27C1,
32'hBED8085B,
32'hBF8D5258,
32'h3EE4C66C,
32'h3E7A9E4E,
32'h3F7D4799,
32'hBD5CE8F2,
32'hBE9294B4,
32'h3F058732,
32'hBEEEA4AF,
32'h3EB99C05,
32'h3C0116CD,
32'h3F14238F,
32'h3E72D197,
32'h3DFBAE29,
32'hBF5BED43,
32'h3E664CCF,
32'hBEE51573,
32'hBF3694FF,
32'h3E9A1FBF,
32'h3E81E453,
32'h3E31C8FC,
32'hBD1A075E,
32'h3C687A64,
32'hBF4DC122,
32'hBE414DA5,
32'hBF7C1B90,
32'hBE20CD24,
32'hBEA64B91,
32'hBF41C6D5,
32'h3E954202,
32'hBE88DA55,
32'hBF8F2FC3,
32'hBCB3D710,
32'h3E2611ED,
32'h3E8922B9,
32'h3E16C67B,
32'h3E8EA388,
32'hBDCF16A4,
32'h3F028ACC,
32'h3F0973F3,
32'hBF53F0C2,
32'h3EDCBAE7,
32'h1DF9D7B2,
32'hBF004096,
32'hBFCAF12E,
32'hBEC8B237,
32'hBF6FA082,
32'h3F070956,
32'h3DAD1D5F,
32'hBED5B03A,
32'hBEE51FC2,
32'hBDA33A61,
32'h3CEB5F51,
32'hBF0EEC78,
32'hBD85CA00,
32'hBF81DBB9,
32'h3E724F1F,
32'hBEDD3186,
32'hBF6781B8,
32'h3E40CC47,
32'hBE7AC610,
32'hBFA10A90,
32'hBE03CE01,
32'h3DADBAB3,
32'h3EFE36AB,
32'hBE7E5FED,
32'h3DE991CC,
32'hBE612230,
32'h3EBE869E,
32'h3F07BE0E,
32'hBF4DC555,
32'h3EBC1AF1,
32'hBE6FEE19,
32'h3DDF1F96,
32'hBFB4BAB1,
32'h3D181DA1,
32'hBF1F72D1,
32'h3F2EB411,
32'h3E198678,
32'hBE8CF13C,
32'hBE13B4A4,
32'hBD801DA7,
32'hBD6EBFA3,
32'hBF31D5F1,
32'hBE1C626C,
32'hBF810A0F,
32'hBE3A1B2E,
32'hBED8F982,
32'hBFA87637,
32'h3E1FFFED,
32'hBF8BFC6C,
32'hBF348B52,
32'hBD2BDF47,
32'h3D272E4A,
32'h3F0D2CAD,
32'h3E4B9E2C,
32'h3F828B13,
32'h3E75F649,
32'h3E600F3D,
32'h3E50033A,
32'hBFC129E8,
32'h3EA2DA77,
32'h3FBDCE1D,
32'h3F30C7E2,
32'h3EA4C46C,
32'hBF9A67D8,
32'h3ECCD456,
32'h3F0EBBFB,
32'h3D64821B,
32'hBE82E867,
32'hBE55DCBC,
32'hBD3D6129,
32'h1DEB9D33,
32'hBE6E4D50,
32'hBE4FFEA4,
32'hBD3F2A4D,
32'hBF21EC6A,
32'h3D365E56,
32'hBF2C1E65,
32'hBD948636,
32'hBF7478BB,
32'hBF8A8027,
32'hBE868AE7,
32'h3DE71960,
32'h3E2FB451,
32'h3CF78F4D,
32'h3F6ADA2E,
32'h3E9FA16D,
32'h3E9DE5B0,
32'hBEB5A690,
32'hC00841F3,
32'hBC5B9E80,
32'hBF07E872,
32'hBDE60620,
32'hBF716C9E,
32'h3EA432B1,
32'h3E0ED793,
32'h3F82BFC6,
32'hBE54D9BD,
32'hBE60902C,
32'hBEFC97AF,
32'hBD708464,
32'hBCDBA1CA,
32'hBE3B366E,
32'hBE209F8C,
32'hBF031504,
32'h3EB8F3BA,
32'hBDFA3A08,
32'hBF603368,
32'h3E2C679E,
32'hBE03C224,
32'hBF9ECDD6,
32'hBE32652A,
32'h0EC1173D,
32'hBE9503FE,
32'hBF029976,
32'hBE61139F,
32'h3EC31DD3,
32'hBEB9C16E,
32'hBF16DF78,
32'hC0076DEA,
32'hBCE051B3,
32'hBE819C50,
32'hBF893658,
32'hBF24C4B0,
32'h3F5C1B08,
32'h3D11DB8A,
32'h3F25329F,
32'h3F5D4F0B,
32'hBF2EA616,
32'hBD24323A,
32'hBD513DCC,
32'hBDC365B9,
32'hBF2E602A,
32'hBDAFA623,
32'hBE48DDF5,
32'h3E887D24,
32'hBDBF287B,
32'hBFB95531,
32'h3F196FF0,
32'hBF2E4B92,
32'hBFD81AC7,
32'h3E9FBCBF,
32'h1DF5D77A,
32'hBF201B4D,
32'hBF318A53,
32'h3DC3AC5F,
32'h3E457606,
32'h3F431A60,
32'hBDA22B33,
32'hBFB1F7BB,
32'h3CAB05F3,
32'h3E829A16,
32'hBEC2F976,
32'h3D93DB11,
32'h3EF097E7,
32'hBD723395,
32'h3F5027F8,
32'h3F597137,
32'hBE5A977D,
32'h3CF1A10A,
32'hBCB1C1E8,
32'hBC132DA6,
32'h3E7B4B66,
32'hBEA59DCF,
32'hBE479ADB,
32'hBF00639B,
32'hBD90FA04,
32'hBF879AEC,
32'hBD284D76,
32'hBF903ABB,
32'hBFD0C0B5,
32'h3F23FE7F,
32'hBCD4E701,
32'hBCB2B056,
32'hBDF1A88F,
32'h3EF9BBC9,
32'h3F128600,
32'h3EA3582A,
32'hBCA2C398,
32'hBF6FF93A,
32'hBDAA8D6A,
32'h3F892F29,
32'h3C9AD739,
32'h3E189064,
32'hBF4E016B,
32'hBDEDD8A7,
32'h1DC9547F,
32'h3F2503EA,
32'h0759A728,
32'hBDA3350D,
32'h3D81ADA0,
32'h3D3847E7,
32'h3E7F2F35,
32'h3C7EE00F,
32'h3DE2B551,
32'h1DCFE0AE,
32'h5DEC7EAD,
32'hBF3BD2B2,
32'h3EFC9EAF,
32'hBE23CE8C,
32'hBF823C52,
32'hBDC5A393,
32'hBD40178C,
32'hBE561E07,
32'hBDA36C26,
32'h3EBE1907,
32'h3F0F7DF4,
32'h3F0F746F,
32'hBD583C9C,
32'hBF248862,
32'h3C777CD8,
32'hBE78EC17,
32'hBC74DE7E,
32'h5DD574DE,
32'h3E868CAD,
32'h1DC0B416,
32'hBCC8A5E6,
32'hBDB01E80,
32'h3DE9C6E6,
32'hBD04D180,
32'hBD38127F,
32'hBDBE0601,
32'h3EA8D967,
32'h3D5F4DBB,
32'hBD261F0A,
32'h3F2A36B7,
32'h3C0937D8,
32'hBD42FB64,
32'h3F233232,
32'h3E92F0B8,
32'h3E242F65,
32'hBEEF3DED,
32'hBCE1551C,
32'hBF1ED5EE,
32'h3DD171F6,
32'hBEC4A37D,
32'hBCA9DB51,
32'h3D1B6AE8,
32'h1DC14AAA,
32'hBE0BF3C8,
32'hBDB821D0,
32'hBDA73BB3,
32'h3D8A4E8C,
32'hBD8AF4D3,
32'h1DF83902,
32'hBE2DDADD,
32'hBDAF3813,
32'hBD4570BF,
32'hBCBE6206,
32'h3C84E289,
32'h0EC1FEB3,
32'hBCAD7034,
32'h3D01183E,
32'hBD236214,
32'hBD03E00E,
32'h3CA6B3D2,
32'h1DEDB196,
32'hBDB44562,
32'h3D90EBFA,
32'hBD7CD23E,
32'h0EDAD526,
32'h3D87E193,
32'h3DA1D895,
32'hBC84658C,
32'hBD6C4914,
32'h3C4A2E7E,
32'h5DCBB534,
32'h3DD4FD0A,
32'h3C1E8A38,
32'hBC307563,
32'h3C3F708F,
32'h3CE99A2A,
32'h3C37799B,
32'hBDEB0AC8,
32'h3D0F1940,
32'hBD09A36C,
32'h3D578126,
32'h3CC00073,
32'h2ECAAE37,
32'h3CB9B2A4,
32'hBA4245F,
32'h3D76DB8D,
32'hBDA8A077,
32'hBCA3E40C,
32'h3D049553,
32'h3CE19E16,
32'hBD1C6B84,
32'hBD1C6239,
32'h3CB59AF5,
32'h3D0A9CFC,
32'hBC2FCED6,
32'hBD8D70C0,
32'hBDD86013,
32'h3D77B9A8,
32'hBD362569,
32'hBD1EACCC,
32'hBD8E6D66,
32'hBCCAEA58,
32'hBD678EAD,
32'h2ECBCEE8,
32'h0EC9133A,
32'h1DD813BE,
32'h3D3C3AD3,
32'h3C09341C,
32'hBCD308F8,
32'hBD32090D,
32'h2E5E28E,
32'hBC2F8EDD,
32'h3D3178D3,
32'h3CE96699,
32'h3D1FFE55,
32'hBC87A4BA,
32'h3D93D986,
32'h3D38ADC9,
32'h3CA09BDB,
32'h5DC84927,
32'h3CAF74E8,
32'hBD38EAD2,
32'h3D95DA73,
32'hBCBBD143,
32'h3C7C3940,
32'hBC5D728D,
32'hBD3D0775,
32'h3D01D96E,
32'hBD66230F,
32'h3C8E0581,
32'hBCC11EA3,
32'h3D106D63,
32'hBD8105DC,
32'hBD65C006,
32'hBD9753D6,
32'h3D846F6D,
32'hBD46FDE7,
32'h3DBFDA3E,
32'h3D287618,
32'h3DCC636B,
32'hBCD64C69,
32'h1DC9AE3D,
32'hBDA42D29,
32'hBCE2A213,
32'hBD1F9023,
32'h3D2092DD,
32'hBDC33104,
32'hBD40EFDB,
32'hBD57E8C5,
32'hBCA8369F,
32'h3D261E67,
32'h3D49F911,
32'h0ED79610,
32'h3CFFBE15,
32'hBD3757D6,
32'h3D36A540,
32'hBCF8831D,
32'h3DB4D64F,
32'hBD849ACC,
32'hBDA96895,
32'hBC12B14A,
32'h3D5BDA24,
32'h5DF63C62,
32'h5DEC3305,
32'h3D497296,
32'hBD393637,
32'hBC2B4F0F,
32'h3DAADD4A,
32'hBCC95DA3,
32'hBD7DFEB4,
32'h3C4083FC,
32'hBC526D59,
32'h3D814FA3,
32'hBDA52275,
32'h3D055AA9,
32'h3D785664,
32'hBD167156,
32'h3D462431,
32'h3CE2AA47,
32'hBC0366FA,
32'h3D4D53F6,
32'hBDE1465A,
32'h3C7F2EB1,
32'h3CC627AC,
32'h3DC2C6D0,
32'h3DDA85CA,
32'h3DDCB456,
32'h3D3A765F,
32'h3D877BE3,
32'h1DF27E07,
32'hBD1E064F,
32'h3DB72938,
32'hBD78FAD5,
32'h3DA59C7F,
32'hBCA2016D,
32'hBD865AED,
32'hBC59193B,
32'hBD39B8C5,
32'hBCCF87FD,
32'hBDE090D0,
32'h3DB1CA6B,
32'h3CA7A364,
32'h3D57B042,
32'h3CD54BE8,
32'h3DCEE565,
32'hBD48D3C6,
32'h3D2AF223,
32'hBDABF5A2,
32'h3CCC2991,
32'hBC9FCB22,
32'hBD84AC84,
32'hBD545A2D,
32'h3DA2B555,
32'h5DE3DDF9,
32'h3C62375B,
32'h3C9F3F05,
32'hBD075EAA,
32'hBC300200,
32'h3D1994FF,
32'hBDA2BD7D,
32'hBCA60176,
32'hBD22F6A3,
32'h2EC65767,
32'h3C6DC94F,
32'hBCFBCEF9,
32'hBDDC1C56,
32'h3DEAE9CC,
32'hBD50CF06,
32'hBDBC3D53,
32'hBCEE1369,
32'h3CDDF873,
32'h3D1946EB,
32'h3D8BF271,
32'hBCAD558B,
32'hBD22C2F5,
32'h3C678DC0,
32'h3C0BE11E,
32'h3D975EC6,
32'h3C8DAC8E,
32'hBD9231B3,
32'hBCE63A94,
32'h3D2FDB34,
32'h3DAE5245,
32'hBD07261D,
32'h5DE25BD9,
32'h3D2742B0,
32'h3D3CD551,
32'h3C73AC8F,
32'h3CD6A33E,
32'hBDCF6D20,
32'hBC998BB6,
32'hBCE02E84,
32'hBD2F61E8,
32'h2E4900E,
32'hBD90BB40,
32'h3D5371CC,
32'h3E06E0B8,
32'h3D599202,
32'h3EDD1947,
32'hBE140F83,
32'h3D3F9852,
32'h3D62CE2B,
32'h3DD4E982,
32'h3C806A42,
32'hBD2FD4F9,
32'h3D09E813,
32'h3D9ED9CB,
32'h3D83FDA4,
32'h3E44FDAF,
32'hBE987FD8,
32'h1DE118B5,
32'hBCD6B307,
32'h3E15A2EE,
32'h3D13A1F3,
32'hBC826CF0,
32'hBE52DEC4,
32'h3D5107E3,
32'hBF3DFF6E,
32'h5DCA42BE,
32'h3F4CB11A,
32'hBE2E9508,
32'h3E9FF273,
32'h3C99B089,
32'hBD784650,
32'hBE2D741B,
32'h3F54CB33,
32'h3E221295,
32'h2ECC69FA,
32'h3F4EEF6F,
32'hBD59488E,
32'hBDDAB86B,
32'hBDC6E6FC,
32'h3DAAB1DD,
32'h3E3F2DDA,
32'h3DB55D31,
32'hBD98F450,
32'hBD1C0E7A,
32'hBD2CFFF5,
32'h3E929A8B,
32'hBF20127E,
32'h3CF08D2F,
32'hBC5ABCFD,
32'h3F37B767,
32'h3EE77C1A,
32'hBE23657F,
32'hBEFCC183,
32'hBDA1DD65,
32'hBF4739A7,
32'h3C284F86,
32'h3F734B71,
32'hBEBF50E5,
32'h3E937D88,
32'hBD9DE9BF,
32'hBE2A3218,
32'h5DF64AD2,
32'h3F1B0ABE,
32'h3DBD4614,
32'hBE7F3645,
32'h3EC2B75A,
32'hBE00E927,
32'hBE854A87,
32'h3CA71840,
32'h3D11A2B3,
32'h3E0CB221,
32'hBDA68FA5,
32'h3DC83B74,
32'hBC4D41BF,
32'hBD99CD53,
32'h3E897E00,
32'hBEBF935B,
32'hBD33C336,
32'hBEC05765,
32'h3E209C11,
32'h3DDAD7E2,
32'hBFAC1326,
32'h3DD12EA2,
32'h3C4F7EB4,
32'hBE8CFEBE,
32'hBDB3DC0C,
32'h3F0B3FB5,
32'h3D179DEA,
32'h3DEF83F4,
32'h3C1E5843,
32'hBF1CBB23,
32'hBCB89075,
32'h3F1B4911,
32'h3E379FF8,
32'hBE11B1DA,
32'h3E4C018B,
32'hBD8B7DE3,
32'hBEE3DE16,
32'hBC2622F6,
32'hBD5FBBFD,
32'h3DE06A7C,
32'hBCBF6D84,
32'h3CC55A95,
32'hBD8D1B4F,
32'hBD5ECA1E,
32'h3E459E2D,
32'hBE80368B,
32'h3D431965,
32'hBED73D90,
32'hBE0A1282,
32'hBE20B1BC,
32'hBFB440C0,
32'h3E469A4F,
32'h3D69197B,
32'h3EAD0F9D,
32'hBD0C2172,
32'h3E409ED7,
32'h3E3F01D3,
32'h3E641017,
32'h3D99C842,
32'hBF392107,
32'hBC555AC8,
32'h3F2E99B1,
32'h3E628299,
32'hBC11B57E,
32'hBE1962B0,
32'h3DBAF50A,
32'hBED2B617,
32'h3D7F877B,
32'hBC8F1DD4,
32'h3EA3CF61,
32'h3CE92DFE,
32'h3C87D61D,
32'h3D264BC8,
32'h3D1654E1,
32'hBD8CD8C8,
32'hBEC15084,
32'hBD18483D,
32'hBEE72708,
32'h3D36FD15,
32'h3E3A307D,
32'hBFB6B2F8,
32'h3DE5E768,
32'hBD90B4F3,
32'h3EBA2F31,
32'hBCA5D5A2,
32'h3E0F5150,
32'h3E6181E4,
32'h3E3921E9,
32'hBC66128D,
32'hBF5994B3,
32'h3F09295D,
32'h3F784EB2,
32'h3F26A6C3,
32'hBE116FAB,
32'hBD99B612,
32'hBCC4106B,
32'h3D19393F,
32'h3EED1EDE,
32'hBE2EE88C,
32'h3EACD4D9,
32'h3C5B0194,
32'h3DD03F15,
32'h3DAE748E,
32'hBDC85832,
32'hBE6A8C3C,
32'h3E5217DD,
32'h1756D033,
32'hBEE79589,
32'h3E6345FE,
32'h3E8DAC83,
32'hBFA69656,
32'hBF4A2899,
32'h5DDA8AFF,
32'hBD9D33A9,
32'hBDD3F0A7,
32'h3E335576,
32'hBE669E46,
32'hBE365B25,
32'h3A44BAE,
32'hBF5E37EB,
32'h3E090C33,
32'h3E169A8D,
32'h3F433EDA,
32'hBDD509ED,
32'h3F0980AB,
32'h3E83AAE1,
32'hBE0FDC22,
32'h3F1713AE,
32'h3D66EF51,
32'h3E85A26F,
32'hBC601334,
32'hBD18CC97,
32'h3DFC3BC2,
32'hBD3161D9,
32'hBE8ECBD1,
32'h3E408637,
32'h3C74FADB,
32'hBE76ED68,
32'h3EC3F7E4,
32'h3D8BE393,
32'hBF61730F,
32'h3E42A36E,
32'h3D838CF1,
32'hBF4ACB3B,
32'hBE784C2A,
32'h3F4B7465,
32'hBDF37C72,
32'hBE70A239,
32'h17504BC7,
32'hBF11D661,
32'h3E07F9EB,
32'hBE8F2F9B,
32'h3F5A06B4,
32'hBE044BB3,
32'h3F430AF2,
32'h3E0A45BD,
32'hBECB6AC8,
32'hBED2A024,
32'hBF24D445,
32'h3E9B3AEB,
32'hBDAC5703,
32'h3C308C14,
32'h3DB28273,
32'hBDF289EF,
32'hBEE527BF,
32'h3E83C181,
32'hBD132FF2,
32'hBED139CD,
32'h3C9DEFE8,
32'hBE06564C,
32'hBF7CF2BA,
32'h3E777B85,
32'h3DA4FEAF,
32'h3E93365D,
32'hBEA95BA7,
32'h3CBFE483,
32'h3CC9E551,
32'hBE816C8C,
32'hBDC1CF29,
32'hBEE45A18,
32'h3DF19E51,
32'h3F12F9B7,
32'h3EE16BF5,
32'h3C40C213,
32'h3E318F36,
32'h3E867CD3,
32'hBE81D6AA,
32'hBD56D3D5,
32'hBF133263,
32'h3ECA9A94,
32'hBD6F2ECF,
32'hBCD04E83,
32'h3E394D77,
32'hBD88B8E3,
32'hBE732B5B,
32'hBEB79B29,
32'h3CC323C8,
32'hBEC6D80E,
32'h3E924FB5,
32'h3F132357,
32'hBF5166B5,
32'h3E01741F,
32'h3CDB5775,
32'h1DC89003,
32'hBEA92B49,
32'h3EF8340E,
32'hBE1DB276,
32'hBDD0FD92,
32'h3CC857E7,
32'hBF41DD96,
32'h3E9D6314,
32'h3EC8A25D,
32'h3EAECDC3,
32'hBE1AACAE,
32'h3ED8E809,
32'h3E653C6D,
32'hBDE1BDAB,
32'h3E642CD8,
32'hBF2865C1,
32'h3E539F58,
32'h1DE87216,
32'h1DC969B0,
32'hBD5A6109,
32'h2ED51635,
32'h3CE0A2AA,
32'hBEB6E030,
32'hBE988844,
32'hBEECA5D0,
32'h3F285C3F,
32'h3F813E35,
32'hBFB6326C,
32'h3EC764CC,
32'hBD83637C,
32'hBDEF0DFB,
32'hBEE88694,
32'h3EAAC66E,
32'hBCEE70D4,
32'h3D356567,
32'hBC51D66E,
32'hBF71568D,
32'h3F2775A5,
32'h3ED0EA77,
32'h3E4FA22B,
32'hBEA2D649,
32'hBD885711,
32'h3E1CAF55,
32'hBEE61ADF,
32'hBED66352,
32'hBEF8DF28,
32'h3E85E6DF,
32'hBD32A3E0,
32'h1DD765F4,
32'hBE2E1DA4,
32'hBC98B3A7,
32'hBEA24EA7,
32'hBD10F134,
32'hBE1BE99F,
32'hBF04065C,
32'h3F39B5DF,
32'h3F86BE7F,
32'hC00C34CB,
32'h3F459373,
32'h3D818829,
32'hBE0BB924,
32'hBEAE150C,
32'hBEB01506,
32'h3ECD49E9,
32'h3E04C8DE,
32'h3C826D85,
32'hBFD9CB6D,
32'h3DDD0E14,
32'hBE932E92,
32'h3D40E926,
32'hBE71FAF4,
32'hBE6749B0,
32'h3F3B63E9,
32'hBE62030B,
32'hBF5268D1,
32'hBEE25B37,
32'h3E173FE3,
32'h3C851B1B,
32'h3DA6D1D0,
32'hBE0C358E,
32'h3CE7DA75,
32'hBDAC3E92,
32'h3F529AC1,
32'hBD5E4AF0,
32'hBD385620,
32'h3F2C086B,
32'hBEF3B734,
32'hBE28B9BF,
32'h3EE68AF6,
32'h3D8648FE,
32'hBD567851,
32'hBE8A6089,
32'hBF2DAE08,
32'h3F61B8FA,
32'hBE1F3664,
32'hBD63E2DA,
32'hBF220E45,
32'h1DFE0C6E,
32'h3ED3E5B6,
32'h3E0D1248,
32'hBE5FFF76,
32'h3DAE5B0F,
32'hBE4BB84E,
32'h3D7C9BAA,
32'h3E144C81,
32'hBE28BDB9,
32'h3E99C993,
32'hBC8A0E77,
32'hBD93CFE6,
32'hBDD1FEA6,
32'h3D00927B,
32'h3E41F84E,
32'h3F1E5125,
32'hBC34F3D1,
32'hBF10C930,
32'h3E79CDB6,
32'h3F227135,
32'hBF05D4C1,
32'hBD96E9FC,
32'hBDA42E34,
32'hBDB5255D,
32'h3E1D92D8,
32'h3F500003,
32'hBEEA9622,
32'hBDAF2446,
32'h0ED15119,
32'hBDD5B67A,
32'h3E3A6677,
32'h3EF5FA3B,
32'hBE1D4137,
32'h3E955CB8,
32'hBE48ED4D,
32'h3DFCD7AD,
32'hBE7F8C3D,
32'hBE3DE8C8,
32'hBEEA5889,
32'h3EA6FDA1,
32'hBCB8B7BC,
32'h3CCED1DF,
32'hBE0B2A50,
32'h1DC28003,
32'h3F057948,
32'h3E4070CE,
32'hBE13E065,
32'hBF0478CF,
32'h3F83C35C,
32'h3E9E05DB,
32'hBE3CDD85,
32'hBEBC38B8,
32'h3D4CE0EE,
32'hBEA983C9,
32'hBE5DBB76,
32'h3EA6A89A,
32'hBE515B6A,
32'hBEF50CAE,
32'h3DDBA051,
32'hBF6E109F,
32'h3E88E5E3,
32'h3F7DD933,
32'h3D11C661,
32'h3EB52654,
32'hBE6D57DE,
32'hBCA6D9B8,
32'hBEADF757,
32'hBE67855F,
32'hBE796DC9,
32'hBE4A7C93,
32'hBDB8C625,
32'hBD13A857,
32'hBE4BCB45,
32'hBCA069ED,
32'hBE296DCE,
32'hBE41A557,
32'h3C83B8B7,
32'hBE93DA0B,
32'h3F8F748C,
32'hBDF8156C,
32'hBE8552EE,
32'h3CB05976,
32'h3D0ED78E,
32'h3E974568,
32'h3E34D3CF,
32'h3D08514F,
32'hBEA8182E,
32'hBF383B29,
32'h3D59CFAA,
32'hBF6C191E,
32'h3E64B2E9,
32'h3F00431B,
32'h3CF28123,
32'h3EACB22D,
32'hBE58B60C,
32'h3CC4D059,
32'h5DF6FBA3,
32'hBD24F220,
32'hBDF711FE,
32'h3E0CA496,
32'hBC12F3C8,
32'h3C3181B2,
32'hBE07364F,
32'h2EC1846F,
32'h1DEE5F7D,
32'hBE45A9B0,
32'hBDE68564,
32'hBECDC65A,
32'h3DB5842F,
32'hBE40BF63,
32'hBF43022F,
32'hBDEAA87F,
32'h3D739AAC,
32'h3ED893AF,
32'hBF3BC62B,
32'hBCC1903F,
32'h3EA87531,
32'h3ECABDD1,
32'h3CAF1BFE,
32'hBEDC7355,
32'hBD22E516,
32'h3E219A9D,
32'h3D031589,
32'h3E57CF55,
32'hBD72874D,
32'h3D07B065,
32'h3DFE705F,
32'hBD914CC2,
32'hBE1EDE34,
32'hBDD3215D,
32'h3C29FD7F,
32'h3CBC0F75,
32'hBDF05ED6,
32'h3CE45A8A,
32'hBE503C67,
32'hBCBDBF68,
32'hBD1E9DA3,
32'hBEBF26B7,
32'h3D0974A5,
32'hBE6604AD,
32'hBE147761,
32'hBEDA7AC5,
32'h3D9B8594,
32'h3EDCE0AB,
32'hBF35345D,
32'hBE1BD65D,
32'hBEF8435D,
32'hBDA47183,
32'h5DD0BBEE,
32'h3C1E3C4C,
32'hBD5B67B6,
32'h3F43BD6D,
32'hBE46CC27,
32'h3E32D53F,
32'h3EAB8D4E,
32'h3D5D0B62,
32'h3D97CF94,
32'h3EECFB86,
32'hBE1298D1,
32'hBC734171,
32'h3DB6BDC0,
32'h3D0DC21A,
32'hBF3C28FA,
32'hBC343C97,
32'hBD4B6EC3,
32'hBED621CC,
32'h3DE8FAEC,
32'hBF08ADD1,
32'h3EAB2697,
32'hBD885644,
32'hBF80648F,
32'hBF332A2B,
32'h3D461FA0,
32'hBDD06507,
32'hBEC4C2CE,
32'hBE9785DB,
32'hBF1C7D1B,
32'h3EF06360,
32'h3C102C72,
32'hBE8DDEF2,
32'h3D5A4FE4,
32'h3EDC3965,
32'hBE167F4A,
32'h3D5E4F3C,
32'hBCFB91F4,
32'hBD6FC103,
32'h3C866576,
32'hBD0624A4,
32'hBDE73E5A,
32'hBC88CD4B,
32'h3CF7440B,
32'hBDE5F13A,
32'hBDAAA2F7,
32'h3CA9B456,
32'h3D222465,
32'h3E3C1141,
32'hBD25F95E,
32'h3E9E0A9D,
32'h3E572450,
32'h3E100A0C,
32'hBC3708E9,
32'hBDD5BDFC,
32'hBC039650,
32'hBE77BC96,
32'hBEB96A12,
32'hBE93AA03,
32'hBDBA39D8,
32'h3E2B5CCC,
32'hBCA1C99B,
32'hBDBF2555,
32'h3C9630A5,
32'h3F069D09,
32'hBD46F654,
32'hBC608E68,
32'h3EA4E25B,
32'hBD7302F9,
32'h3D62C50C,
32'h3E4F01CC,
32'h3A1D2D0,
32'h5DF12FE7,
32'hBDC39C14,
32'hBD81488C,
32'h3CCD4CB0,
32'hBD77B855,
32'hBCBE8CF4,
32'hBED215AB,
32'h3D659A87,
32'hBD72C444,
32'h3EB91BB6,
32'h3E0F83EA,
32'hBD97A563,
32'hBE0FED19,
32'h1DF3ECF0,
32'hBEF160F8,
32'h3D6C95C1,
32'h3EC9C6BB,
32'hBD9D8D41,
32'h3EEE45E6,
32'hBC882877,
32'hBECA23DB,
32'hBD78D7A8,
32'h3C641BF7,
32'h3CC57A12,
32'hBC68A478,
32'h5DCA4F3A,
32'h3DD4232E,
32'h3D51AB3A,
32'hBC40BFE1,
32'h3CBEB8F0,
32'h5DF8C42F,
32'h3C2B6009,
32'hBC0A3779,
32'hBD5795B1,
32'hBDC095E0,
32'h3D8BFF6F,
32'hBD80C4FD,
32'h2EDDCA53,
32'hBD105FB6,
32'hBCF3E922,
32'hBD598BA5,
32'h3D8A86AE,
32'h3C596503,
32'hBCE883EF,
32'h3D256831,
32'h3DC427D1,
32'h3DCC5257,
32'hBD2FF0AA,
32'h1DD5EC77,
32'h3D26AB58,
32'h0EDE7301,
32'hBD2DAA9A,
32'hBD56CBF2,
32'h3DDC0B42,
32'hBD397AC9,
32'h3C0601AD,
32'hBCFAB8E6,
32'hBD868B68,
32'hBD8FE5CD,
32'h1DED207A,
32'h3CF6A362,
32'h3D9235BE,
32'hBD1FEA15,
32'h3D163005,
32'h3D1EC23A,
32'hBC5CB342,
32'h0E58517,
32'hBD00F8DA,
32'hBD39B723,
32'h3D1FB638,
32'hBD2F09FB,
32'hBDE46AA8,
32'h5DE883DE,
32'h5DC2089B,
32'hBCE9296E,
32'h3DE61BEE,
32'hBD0B1369,
32'h3DB3C020,
32'hBCA0986D,
32'h3D7D50D9,
32'hBD198006,
32'h3D93B673,
32'h175DFD59,
32'hBC5FDCAA,
32'h3D31E46C,
32'hBD3C0F6A,
32'h3D0CCC60,
32'h3D9ADFB6,
32'hBD312B6C,
32'hBD7120F4,
32'h2ED0ABA6,
32'h3D3DAEA3,
32'h3DAB0088,
32'hBD735ABA,
32'h3D667F7B,
32'hBD659DB5,
32'hBD642380,
32'h3C3900DC,
32'h3C9DE3D2,
32'h3D945B31,
32'h5DD915EC,
32'hBDE830DD,
32'h3CB4498F,
32'hBD9381E0,
32'hBD37BB4F,
32'hBCAB328F,
32'h3D6431C1,
32'h3D1E6E46,
32'h1DF91C02,
32'hBD84C236,
32'h3D23543A,
32'hBD9C86E1,
32'h3D7C6FAE,
32'h1DCF9DD7,
32'hBD900EBB,
32'hBA35559,
32'hBD43CB2F,
32'hBCD13634,
32'hBD0FC1E2,
32'h3DD9F273,
32'hBDAD5BC1,
32'hBC3D1EE8,
32'hBD01D747,
32'h3D7C3991,
32'hBC66514A,
32'hBD5CE8D5,
32'h3CC768FF,
32'h3D49FDE7,
32'hBD57966A,
32'hBD202830,
32'hBD56CE81,
32'h3CA0A169,
32'hBD4C40C4,
32'hBCF2FF73,
32'hBC6BCB48,
32'hBDD52812,
32'h3D462B0F,
32'hBC802175,
32'h3DDAF18B,
32'hBD9445A5,
32'hBDAD16D3
};

	assign weight = ROM[addr];

endmodule 