module memory_parser;

parameter size = 47040;

task memory_contents(output logic[15:0] mem_array[0:size-1]);

mem_array[1] = 16'hc54c;
mem_array[0] = 16'hbcd6;
mem_array[3] = 16'h1706;
mem_array[2] = 16'h3d82;
mem_array[5] = 16'h7bf2;
mem_array[4] = 16'h3d31;
mem_array[7] = 16'h0db5;
mem_array[6] = 16'hbcdd;
mem_array[9] = 16'hd9f1;
mem_array[8] = 16'hbd88;
mem_array[11] = 16'h3af5;
mem_array[10] = 16'hbc46;
mem_array[13] = 16'h508c;
mem_array[12] = 16'hbd1e;
mem_array[15] = 16'hac22;
mem_array[14] = 16'hbc22;
mem_array[17] = 16'h8956;
mem_array[16] = 16'hbd46;
mem_array[19] = 16'h7352;
mem_array[18] = 16'hbd7d;
mem_array[21] = 16'h0974;
mem_array[20] = 16'hbc7f;
mem_array[23] = 16'h1565;
mem_array[22] = 16'h3d63;
mem_array[25] = 16'ha41a;
mem_array[24] = 16'h3d97;
mem_array[27] = 16'h33cc;
mem_array[26] = 16'hbd4e;
mem_array[29] = 16'h3006;
mem_array[28] = 16'hbd83;
mem_array[31] = 16'h4a1d;
mem_array[30] = 16'h3ce9;
mem_array[33] = 16'h80de;
mem_array[32] = 16'hbd01;
mem_array[35] = 16'h8610;
mem_array[34] = 16'hbd3b;
mem_array[37] = 16'h378e;
mem_array[36] = 16'hbd19;
mem_array[39] = 16'h5fc3;
mem_array[38] = 16'h3c7c;
mem_array[41] = 16'h8c5a;
mem_array[40] = 16'h3ca5;
mem_array[43] = 16'h4833;
mem_array[42] = 16'hbd1f;
mem_array[45] = 16'hbf1f;
mem_array[44] = 16'h3d03;
mem_array[47] = 16'h6ea0;
mem_array[46] = 16'hbb7d;
mem_array[49] = 16'hd1b1;
mem_array[48] = 16'h3c8c;
mem_array[51] = 16'h7a36;
mem_array[50] = 16'hbd9d;
mem_array[53] = 16'h2247;
mem_array[52] = 16'h3ce3;
mem_array[55] = 16'h476b;
mem_array[54] = 16'hbd85;
mem_array[57] = 16'h7ea0;
mem_array[56] = 16'hbc13;
mem_array[59] = 16'h2f07;
mem_array[58] = 16'hbc2c;
mem_array[61] = 16'h5e25;
mem_array[60] = 16'h3b58;
mem_array[63] = 16'hec07;
mem_array[62] = 16'h3cd1;
mem_array[65] = 16'h8ff9;
mem_array[64] = 16'hbc0f;
mem_array[67] = 16'ha11e;
mem_array[66] = 16'h3d53;
mem_array[69] = 16'h90ed;
mem_array[68] = 16'h3d15;
mem_array[71] = 16'h1b34;
mem_array[70] = 16'h3d54;
mem_array[73] = 16'heec4;
mem_array[72] = 16'hbd9a;
mem_array[75] = 16'h893a;
mem_array[74] = 16'hbd9a;
mem_array[77] = 16'h29c0;
mem_array[76] = 16'hbade;
mem_array[79] = 16'hbe02;
mem_array[78] = 16'hbd51;
mem_array[81] = 16'h52e7;
mem_array[80] = 16'h3bf0;
mem_array[83] = 16'h2158;
mem_array[82] = 16'hbdb4;
mem_array[85] = 16'hfecf;
mem_array[84] = 16'h3d9b;
mem_array[87] = 16'h9868;
mem_array[86] = 16'h3cff;
mem_array[89] = 16'h8036;
mem_array[88] = 16'h3dba;
mem_array[91] = 16'h6f44;
mem_array[90] = 16'hbca0;
mem_array[93] = 16'h0bb9;
mem_array[92] = 16'h3dc2;
mem_array[95] = 16'hf580;
mem_array[94] = 16'h3ca1;
mem_array[97] = 16'h5644;
mem_array[96] = 16'hbd6a;
mem_array[99] = 16'hcc8d;
mem_array[98] = 16'h3bb8;
mem_array[101] = 16'h25f1;
mem_array[100] = 16'hbd98;
mem_array[103] = 16'h9974;
mem_array[102] = 16'hbcfd;
mem_array[105] = 16'h83a8;
mem_array[104] = 16'hbca7;
mem_array[107] = 16'h360d;
mem_array[106] = 16'hbd2d;
mem_array[109] = 16'ha97b;
mem_array[108] = 16'h3d84;
mem_array[111] = 16'ha216;
mem_array[110] = 16'hbcd2;
mem_array[113] = 16'h45da;
mem_array[112] = 16'h3cbf;
mem_array[115] = 16'h6a1d;
mem_array[114] = 16'hbce3;
mem_array[117] = 16'h94ac;
mem_array[116] = 16'hbd1b;
mem_array[119] = 16'hb4cc;
mem_array[118] = 16'hbcd4;
mem_array[121] = 16'hcf72;
mem_array[120] = 16'h3dbe;
mem_array[123] = 16'hfb28;
mem_array[122] = 16'hbcca;
mem_array[125] = 16'hfab0;
mem_array[124] = 16'hbd30;
mem_array[127] = 16'ha312;
mem_array[126] = 16'h3c85;
mem_array[129] = 16'ha0d4;
mem_array[128] = 16'h3d75;
mem_array[131] = 16'h1df7;
mem_array[130] = 16'h3cff;
mem_array[133] = 16'h849b;
mem_array[132] = 16'hbd8f;
mem_array[135] = 16'h40ca;
mem_array[134] = 16'hbca1;
mem_array[137] = 16'h5eaf;
mem_array[136] = 16'h3c8c;
mem_array[139] = 16'habc4;
mem_array[138] = 16'hbd97;
mem_array[141] = 16'h73a0;
mem_array[140] = 16'hbce6;
mem_array[143] = 16'hf725;
mem_array[142] = 16'h3d4a;
mem_array[145] = 16'hdbf3;
mem_array[144] = 16'h3c85;
mem_array[147] = 16'h29f7;
mem_array[146] = 16'h3db5;
mem_array[149] = 16'h2030;
mem_array[148] = 16'h3d9a;
mem_array[151] = 16'hf1e5;
mem_array[150] = 16'hbce8;
mem_array[153] = 16'h11c7;
mem_array[152] = 16'h3d2c;
mem_array[155] = 16'hf4bd;
mem_array[154] = 16'hbc27;
mem_array[157] = 16'h0244;
mem_array[156] = 16'hbc9a;
mem_array[159] = 16'h49ed;
mem_array[158] = 16'h3de0;
mem_array[161] = 16'ha6cf;
mem_array[160] = 16'hbc3c;
mem_array[163] = 16'hac79;
mem_array[162] = 16'hbd98;
mem_array[165] = 16'h4ae2;
mem_array[164] = 16'h3d1a;
mem_array[167] = 16'hc7e2;
mem_array[166] = 16'hbce8;
mem_array[169] = 16'he4f4;
mem_array[168] = 16'h3c71;
mem_array[171] = 16'h17a1;
mem_array[170] = 16'h3d74;
mem_array[173] = 16'h3ade;
mem_array[172] = 16'hbd58;
mem_array[175] = 16'hf2a6;
mem_array[174] = 16'h3d77;
mem_array[177] = 16'hce9a;
mem_array[176] = 16'h3ca7;
mem_array[179] = 16'hc21d;
mem_array[178] = 16'h3d09;
mem_array[181] = 16'hd628;
mem_array[180] = 16'h3d65;
mem_array[183] = 16'h954f;
mem_array[182] = 16'hbc9c;
mem_array[185] = 16'hf2b1;
mem_array[184] = 16'h3d17;
mem_array[187] = 16'h79f6;
mem_array[186] = 16'hbbc5;
mem_array[189] = 16'h6cdd;
mem_array[188] = 16'hbd39;
mem_array[191] = 16'hfddd;
mem_array[190] = 16'h3d32;
mem_array[193] = 16'h7080;
mem_array[192] = 16'hbdd0;
mem_array[195] = 16'h9cb0;
mem_array[194] = 16'h3db9;
mem_array[197] = 16'h4155;
mem_array[196] = 16'h3c82;
mem_array[199] = 16'hc993;
mem_array[198] = 16'hbd90;
mem_array[201] = 16'hb07a;
mem_array[200] = 16'h3d33;
mem_array[203] = 16'hf1f2;
mem_array[202] = 16'hbdbb;
mem_array[205] = 16'h9691;
mem_array[204] = 16'hbc2e;
mem_array[207] = 16'h5dcb;
mem_array[206] = 16'hbd7b;
mem_array[209] = 16'ha511;
mem_array[208] = 16'hbd0d;
mem_array[211] = 16'h553a;
mem_array[210] = 16'h3ccf;
mem_array[213] = 16'h241b;
mem_array[212] = 16'hbd7c;
mem_array[215] = 16'h7dac;
mem_array[214] = 16'hbd83;
mem_array[217] = 16'hc066;
mem_array[216] = 16'h3db9;
mem_array[219] = 16'hba45;
mem_array[218] = 16'hbd1f;
mem_array[221] = 16'hd1cc;
mem_array[220] = 16'h3ca4;
mem_array[223] = 16'h6f00;
mem_array[222] = 16'hbc81;
mem_array[225] = 16'hcf4f;
mem_array[224] = 16'hbc21;
mem_array[227] = 16'hba0b;
mem_array[226] = 16'h3d64;
mem_array[229] = 16'h7d50;
mem_array[228] = 16'h3d17;
mem_array[231] = 16'h3e96;
mem_array[230] = 16'hbdad;
mem_array[233] = 16'h3918;
mem_array[232] = 16'h3d1e;
mem_array[235] = 16'h7b6d;
mem_array[234] = 16'h3d61;
mem_array[237] = 16'hda78;
mem_array[236] = 16'h3d7f;
mem_array[239] = 16'h8f17;
mem_array[238] = 16'h3d60;
mem_array[241] = 16'h714f;
mem_array[240] = 16'hbc9c;
mem_array[243] = 16'h4a7e;
mem_array[242] = 16'h3d64;
mem_array[245] = 16'h2cda;
mem_array[244] = 16'h3d7f;
mem_array[247] = 16'h5d65;
mem_array[246] = 16'h3cc3;
mem_array[249] = 16'hda2a;
mem_array[248] = 16'h3c99;
mem_array[251] = 16'h717c;
mem_array[250] = 16'hbd19;
mem_array[253] = 16'h31ad;
mem_array[252] = 16'h3c84;
mem_array[255] = 16'h5f51;
mem_array[254] = 16'h3ae5;
mem_array[257] = 16'hd8dc;
mem_array[256] = 16'hbd98;
mem_array[259] = 16'h207a;
mem_array[258] = 16'hbc54;
mem_array[261] = 16'hcf50;
mem_array[260] = 16'hbcb5;
mem_array[263] = 16'h8193;
mem_array[262] = 16'hbdac;
mem_array[265] = 16'h86e1;
mem_array[264] = 16'hbd94;
mem_array[267] = 16'hf692;
mem_array[266] = 16'hbd09;
mem_array[269] = 16'h64db;
mem_array[268] = 16'hbc9d;
mem_array[271] = 16'hc91c;
mem_array[270] = 16'h3b98;
mem_array[273] = 16'h2c64;
mem_array[272] = 16'hbd41;
mem_array[275] = 16'he416;
mem_array[274] = 16'h3cbd;
mem_array[277] = 16'he87c;
mem_array[276] = 16'h3d06;
mem_array[279] = 16'h1b49;
mem_array[278] = 16'h3dbe;
mem_array[281] = 16'h9ec3;
mem_array[280] = 16'h3b95;
mem_array[283] = 16'h535d;
mem_array[282] = 16'h3c7b;
mem_array[285] = 16'h60b9;
mem_array[284] = 16'h3d27;
mem_array[287] = 16'h11a9;
mem_array[286] = 16'h3d12;
mem_array[289] = 16'ha23f;
mem_array[288] = 16'hbbe2;
mem_array[291] = 16'h89b2;
mem_array[290] = 16'hbdb9;
mem_array[293] = 16'hb3bb;
mem_array[292] = 16'hbd27;
mem_array[295] = 16'hf2eb;
mem_array[294] = 16'h3cf5;
mem_array[297] = 16'h2545;
mem_array[296] = 16'hbd1b;
mem_array[299] = 16'h9af2;
mem_array[298] = 16'h3d5f;
mem_array[301] = 16'h1115;
mem_array[300] = 16'hbd88;
mem_array[303] = 16'h435b;
mem_array[302] = 16'h3cbd;
mem_array[305] = 16'h5691;
mem_array[304] = 16'hbcbe;
mem_array[307] = 16'h23cb;
mem_array[306] = 16'h3c00;
mem_array[309] = 16'hab48;
mem_array[308] = 16'h3d71;
mem_array[311] = 16'hf53a;
mem_array[310] = 16'h3d6e;
mem_array[313] = 16'h8619;
mem_array[312] = 16'h3b20;
mem_array[315] = 16'h30b0;
mem_array[314] = 16'hbd75;
mem_array[317] = 16'h41f1;
mem_array[316] = 16'hbcca;
mem_array[319] = 16'he122;
mem_array[318] = 16'hbd92;
mem_array[321] = 16'h0993;
mem_array[320] = 16'hbd8d;
mem_array[323] = 16'h7da9;
mem_array[322] = 16'hbd2f;
mem_array[325] = 16'h1043;
mem_array[324] = 16'h3d8e;
mem_array[327] = 16'h732e;
mem_array[326] = 16'hbd66;
mem_array[329] = 16'h3955;
mem_array[328] = 16'h3d49;
mem_array[331] = 16'h62dd;
mem_array[330] = 16'hbd38;
mem_array[333] = 16'h4c9a;
mem_array[332] = 16'hbd10;
mem_array[335] = 16'hfcaf;
mem_array[334] = 16'h3cc7;
mem_array[337] = 16'hef08;
mem_array[336] = 16'h3c5c;
mem_array[339] = 16'h1226;
mem_array[338] = 16'h3c3d;
mem_array[341] = 16'hb1f6;
mem_array[340] = 16'h3c80;
mem_array[343] = 16'h99b4;
mem_array[342] = 16'hbdcb;
mem_array[345] = 16'h5476;
mem_array[344] = 16'hbc89;
mem_array[347] = 16'ha559;
mem_array[346] = 16'hbd51;
mem_array[349] = 16'hef65;
mem_array[348] = 16'h3cf8;
mem_array[351] = 16'h9847;
mem_array[350] = 16'h3c6e;
mem_array[353] = 16'h3bc3;
mem_array[352] = 16'h3c5c;
mem_array[355] = 16'h8965;
mem_array[354] = 16'hbb8b;
mem_array[357] = 16'he19c;
mem_array[356] = 16'hbc65;
mem_array[359] = 16'hff00;
mem_array[358] = 16'hbd9a;
mem_array[361] = 16'h0b62;
mem_array[360] = 16'hbd77;
mem_array[363] = 16'h6b73;
mem_array[362] = 16'h3bf2;
mem_array[365] = 16'h9e58;
mem_array[364] = 16'hbd42;
mem_array[367] = 16'hba3e;
mem_array[366] = 16'hbb8b;
mem_array[369] = 16'haa89;
mem_array[368] = 16'h3bdb;
mem_array[371] = 16'he5ea;
mem_array[370] = 16'hbcc4;
mem_array[373] = 16'h3c1c;
mem_array[372] = 16'h3d2f;
mem_array[375] = 16'h293f;
mem_array[374] = 16'hbb58;
mem_array[377] = 16'hcc97;
mem_array[376] = 16'hbd98;
mem_array[379] = 16'hab27;
mem_array[378] = 16'h3b83;
mem_array[381] = 16'hb48b;
mem_array[380] = 16'h3b95;
mem_array[383] = 16'ha073;
mem_array[382] = 16'hbd33;
mem_array[385] = 16'haa27;
mem_array[384] = 16'hbd88;
mem_array[387] = 16'h6118;
mem_array[386] = 16'hbacc;
mem_array[389] = 16'hcce1;
mem_array[388] = 16'hbbd3;
mem_array[391] = 16'h39bd;
mem_array[390] = 16'h3c82;
mem_array[393] = 16'h057c;
mem_array[392] = 16'h3cd2;
mem_array[395] = 16'h8eb4;
mem_array[394] = 16'hbcb1;
mem_array[397] = 16'h0dd9;
mem_array[396] = 16'hbb3b;
mem_array[399] = 16'hefe9;
mem_array[398] = 16'h3dc6;
mem_array[401] = 16'h2b97;
mem_array[400] = 16'h3d28;
mem_array[403] = 16'hf3e9;
mem_array[402] = 16'h3d66;
mem_array[405] = 16'h9310;
mem_array[404] = 16'hbc3b;
mem_array[407] = 16'h5f88;
mem_array[406] = 16'hbd24;
mem_array[409] = 16'h0da3;
mem_array[408] = 16'h3d53;
mem_array[411] = 16'hb363;
mem_array[410] = 16'hbcbd;
mem_array[413] = 16'h3bb8;
mem_array[412] = 16'h3d97;
mem_array[415] = 16'h1341;
mem_array[414] = 16'hbcf5;
mem_array[417] = 16'h6071;
mem_array[416] = 16'h3b2d;
mem_array[419] = 16'h3505;
mem_array[418] = 16'hbda8;
mem_array[421] = 16'h891b;
mem_array[420] = 16'hbd70;
mem_array[423] = 16'hb015;
mem_array[422] = 16'h3db0;
mem_array[425] = 16'hdff9;
mem_array[424] = 16'h3d25;
mem_array[427] = 16'h6ee0;
mem_array[426] = 16'h3dce;
mem_array[429] = 16'ha258;
mem_array[428] = 16'h3c98;
mem_array[431] = 16'hccd5;
mem_array[430] = 16'hbc23;
mem_array[433] = 16'h1cc8;
mem_array[432] = 16'hba1a;
mem_array[435] = 16'h6e5a;
mem_array[434] = 16'hbd18;
mem_array[437] = 16'h7135;
mem_array[436] = 16'hbcb0;
mem_array[439] = 16'h9e08;
mem_array[438] = 16'h3d83;
mem_array[441] = 16'h0136;
mem_array[440] = 16'h3d77;
mem_array[443] = 16'h8a8a;
mem_array[442] = 16'h3c2a;
mem_array[445] = 16'h69b9;
mem_array[444] = 16'hbda4;
mem_array[447] = 16'h87f6;
mem_array[446] = 16'h3d11;
mem_array[449] = 16'h5147;
mem_array[448] = 16'h3d9e;
mem_array[451] = 16'h82f1;
mem_array[450] = 16'hbd68;
mem_array[453] = 16'h1600;
mem_array[452] = 16'h3d2c;
mem_array[455] = 16'hfc02;
mem_array[454] = 16'hbdb3;
mem_array[457] = 16'he1e1;
mem_array[456] = 16'h3d33;
mem_array[459] = 16'h50a2;
mem_array[458] = 16'h3c81;
mem_array[461] = 16'h43b1;
mem_array[460] = 16'hbd88;
mem_array[463] = 16'h90c5;
mem_array[462] = 16'h3d38;
mem_array[465] = 16'h9cce;
mem_array[464] = 16'h3d3d;
mem_array[467] = 16'h432e;
mem_array[466] = 16'h3d52;
mem_array[469] = 16'hc99c;
mem_array[468] = 16'hbc63;
mem_array[471] = 16'h7a31;
mem_array[470] = 16'hbbc9;
mem_array[473] = 16'hbb6a;
mem_array[472] = 16'h3d03;
mem_array[475] = 16'ha2d2;
mem_array[474] = 16'h3cfd;
mem_array[477] = 16'h8786;
mem_array[476] = 16'hbc5a;
mem_array[479] = 16'hd034;
mem_array[478] = 16'h3d71;
mem_array[481] = 16'h694e;
mem_array[480] = 16'h3d00;
mem_array[483] = 16'hc885;
mem_array[482] = 16'h3cb0;
mem_array[485] = 16'h3154;
mem_array[484] = 16'hbd9c;
mem_array[487] = 16'ha0d3;
mem_array[486] = 16'h3d89;
mem_array[489] = 16'h3d72;
mem_array[488] = 16'h3d27;
mem_array[491] = 16'hfd4c;
mem_array[490] = 16'h3c14;
mem_array[493] = 16'h8900;
mem_array[492] = 16'h3d5f;
mem_array[495] = 16'hc7b3;
mem_array[494] = 16'hbc21;
mem_array[497] = 16'hf40e;
mem_array[496] = 16'hbc88;
mem_array[499] = 16'h3773;
mem_array[498] = 16'h3cb6;
mem_array[501] = 16'h4116;
mem_array[500] = 16'h3d0b;
mem_array[503] = 16'hd4e5;
mem_array[502] = 16'h3d44;
mem_array[505] = 16'h634e;
mem_array[504] = 16'h3d6a;
mem_array[507] = 16'hc020;
mem_array[506] = 16'hbd03;
mem_array[509] = 16'h6144;
mem_array[508] = 16'hbdd9;
mem_array[511] = 16'h23ac;
mem_array[510] = 16'h3d92;
mem_array[513] = 16'h18d6;
mem_array[512] = 16'h3db4;
mem_array[515] = 16'he39e;
mem_array[514] = 16'h3d5a;
mem_array[517] = 16'h0c6a;
mem_array[516] = 16'hbcda;
mem_array[519] = 16'h07b7;
mem_array[518] = 16'hbc4c;
mem_array[521] = 16'h3614;
mem_array[520] = 16'hbcab;
mem_array[523] = 16'hc439;
mem_array[522] = 16'h3c14;
mem_array[525] = 16'hfcc3;
mem_array[524] = 16'h3c8f;
mem_array[527] = 16'he3ce;
mem_array[526] = 16'hbd38;
mem_array[529] = 16'hb8f3;
mem_array[528] = 16'hbbeb;
mem_array[531] = 16'hed9e;
mem_array[530] = 16'hbcb6;
mem_array[533] = 16'h77e5;
mem_array[532] = 16'hbba8;
mem_array[535] = 16'h81b3;
mem_array[534] = 16'h3dad;
mem_array[537] = 16'h5acb;
mem_array[536] = 16'h3d9e;
mem_array[539] = 16'h5861;
mem_array[538] = 16'h3d4c;
mem_array[541] = 16'h6fda;
mem_array[540] = 16'h3c8c;
mem_array[543] = 16'h0d95;
mem_array[542] = 16'h3d89;
mem_array[545] = 16'ha8cd;
mem_array[544] = 16'hbbb9;
mem_array[547] = 16'ha3ab;
mem_array[546] = 16'hbd02;
mem_array[549] = 16'h0dbf;
mem_array[548] = 16'hbd01;
mem_array[551] = 16'h5a34;
mem_array[550] = 16'h3cae;
mem_array[553] = 16'h3ab0;
mem_array[552] = 16'hbcc2;
mem_array[555] = 16'h9b2b;
mem_array[554] = 16'h3c2e;
mem_array[557] = 16'h9446;
mem_array[556] = 16'h3d92;
mem_array[559] = 16'hdd81;
mem_array[558] = 16'h3da2;
mem_array[561] = 16'ha91f;
mem_array[560] = 16'h3d31;
mem_array[563] = 16'hb720;
mem_array[562] = 16'h3d14;
mem_array[565] = 16'heb78;
mem_array[564] = 16'h3d2e;
mem_array[567] = 16'h95d6;
mem_array[566] = 16'hbd8c;
mem_array[569] = 16'hacfe;
mem_array[568] = 16'h3c97;
mem_array[571] = 16'ha9d7;
mem_array[570] = 16'h3d89;
mem_array[573] = 16'hdb39;
mem_array[572] = 16'hbc62;
mem_array[575] = 16'h7e93;
mem_array[574] = 16'h3d57;
mem_array[577] = 16'hd837;
mem_array[576] = 16'hbcb3;
mem_array[579] = 16'h3124;
mem_array[578] = 16'hb93b;
mem_array[581] = 16'h2f28;
mem_array[580] = 16'hbd10;
mem_array[583] = 16'h54f4;
mem_array[582] = 16'h3cce;
mem_array[585] = 16'ha9ac;
mem_array[584] = 16'h3de9;
mem_array[587] = 16'hf741;
mem_array[586] = 16'h3d0e;
mem_array[589] = 16'he454;
mem_array[588] = 16'hbce2;
mem_array[591] = 16'h83ef;
mem_array[590] = 16'h3d5e;
mem_array[593] = 16'h5399;
mem_array[592] = 16'h3be3;
mem_array[595] = 16'hcbed;
mem_array[594] = 16'hbc62;
mem_array[597] = 16'hf5d0;
mem_array[596] = 16'h3ac6;
mem_array[599] = 16'he555;
mem_array[598] = 16'hbdac;
mem_array[601] = 16'h7538;
mem_array[600] = 16'hbc70;
mem_array[603] = 16'h84c8;
mem_array[602] = 16'h3c86;
mem_array[605] = 16'h6886;
mem_array[604] = 16'h3d48;
mem_array[607] = 16'h6594;
mem_array[606] = 16'hbd3f;
mem_array[609] = 16'h979c;
mem_array[608] = 16'h3d50;
mem_array[611] = 16'hdb26;
mem_array[610] = 16'h3d12;
mem_array[613] = 16'he718;
mem_array[612] = 16'hbd96;
mem_array[615] = 16'hde34;
mem_array[614] = 16'h3d37;
mem_array[617] = 16'h2a3c;
mem_array[616] = 16'h3d1b;
mem_array[619] = 16'h56b6;
mem_array[618] = 16'hbd37;
mem_array[621] = 16'he987;
mem_array[620] = 16'hbcad;
mem_array[623] = 16'h5b60;
mem_array[622] = 16'h3d57;
mem_array[625] = 16'h59d6;
mem_array[624] = 16'hbdaf;
mem_array[627] = 16'h5c3f;
mem_array[626] = 16'h3d6e;
mem_array[629] = 16'heee9;
mem_array[628] = 16'h3dcc;
mem_array[631] = 16'hc268;
mem_array[630] = 16'h3cf4;
mem_array[633] = 16'he6fe;
mem_array[632] = 16'hbd4f;
mem_array[635] = 16'hdf8f;
mem_array[634] = 16'hbd84;
mem_array[637] = 16'hd9f3;
mem_array[636] = 16'h3cb9;
mem_array[639] = 16'h34a4;
mem_array[638] = 16'hbd2b;
mem_array[641] = 16'h27a7;
mem_array[640] = 16'hbd49;
mem_array[643] = 16'h04c9;
mem_array[642] = 16'hbc9d;
mem_array[645] = 16'h1579;
mem_array[644] = 16'h3c9a;
mem_array[647] = 16'hd9a7;
mem_array[646] = 16'hbb39;
mem_array[649] = 16'he2d9;
mem_array[648] = 16'h3b88;
mem_array[651] = 16'hd566;
mem_array[650] = 16'h3c93;
mem_array[653] = 16'hd878;
mem_array[652] = 16'hbc9e;
mem_array[655] = 16'h4571;
mem_array[654] = 16'h3d07;
mem_array[657] = 16'h59c4;
mem_array[656] = 16'hbdb2;
mem_array[659] = 16'h56fd;
mem_array[658] = 16'hbd08;
mem_array[661] = 16'h0b68;
mem_array[660] = 16'hbbea;
mem_array[663] = 16'h65f8;
mem_array[662] = 16'hbc6c;
mem_array[665] = 16'h8510;
mem_array[664] = 16'hbd22;
mem_array[667] = 16'he635;
mem_array[666] = 16'h3c14;
mem_array[669] = 16'hbcf0;
mem_array[668] = 16'h3d4e;
mem_array[671] = 16'hdf21;
mem_array[670] = 16'hbc0d;
mem_array[673] = 16'hf551;
mem_array[672] = 16'hbcf5;
mem_array[675] = 16'h93f7;
mem_array[674] = 16'h3c1d;
mem_array[677] = 16'h6678;
mem_array[676] = 16'h3db5;
mem_array[679] = 16'h19ef;
mem_array[678] = 16'hbbf9;
mem_array[681] = 16'h5bcb;
mem_array[680] = 16'hbdda;
mem_array[683] = 16'hc61d;
mem_array[682] = 16'h3d7e;
mem_array[685] = 16'h9994;
mem_array[684] = 16'hbd08;
mem_array[687] = 16'hecea;
mem_array[686] = 16'hbda7;
mem_array[689] = 16'h0954;
mem_array[688] = 16'hbcb0;
mem_array[691] = 16'hbd6d;
mem_array[690] = 16'hbc8a;
mem_array[693] = 16'h2c3a;
mem_array[692] = 16'hbd8b;
mem_array[695] = 16'h321c;
mem_array[694] = 16'h3d1c;
mem_array[697] = 16'hac2a;
mem_array[696] = 16'h3d02;
mem_array[699] = 16'h6a8d;
mem_array[698] = 16'h3d93;
mem_array[701] = 16'h2a06;
mem_array[700] = 16'h3c96;
mem_array[703] = 16'h9ddb;
mem_array[702] = 16'h3d13;
mem_array[705] = 16'hba55;
mem_array[704] = 16'hbcc3;
mem_array[707] = 16'h4e59;
mem_array[706] = 16'hbd0f;
mem_array[709] = 16'h1c6f;
mem_array[708] = 16'hbd2d;
mem_array[711] = 16'hc6a1;
mem_array[710] = 16'hbdae;
mem_array[713] = 16'hdfe9;
mem_array[712] = 16'hbbf6;
mem_array[715] = 16'h6b16;
mem_array[714] = 16'hbc05;
mem_array[717] = 16'h9a26;
mem_array[716] = 16'h3dd9;
mem_array[719] = 16'h9e05;
mem_array[718] = 16'hbd8e;
mem_array[721] = 16'h7a76;
mem_array[720] = 16'hbdb5;
mem_array[723] = 16'h0f3c;
mem_array[722] = 16'hbb1d;
mem_array[725] = 16'h355b;
mem_array[724] = 16'h3c94;
mem_array[727] = 16'h8c4f;
mem_array[726] = 16'hbdab;
mem_array[729] = 16'h856b;
mem_array[728] = 16'hbb5d;
mem_array[731] = 16'h8168;
mem_array[730] = 16'h3d46;
mem_array[733] = 16'hff51;
mem_array[732] = 16'h3d8b;
mem_array[735] = 16'h377e;
mem_array[734] = 16'h3d29;
mem_array[737] = 16'h1938;
mem_array[736] = 16'h3a6b;
mem_array[739] = 16'h48c5;
mem_array[738] = 16'h3d8a;
mem_array[741] = 16'hd7fe;
mem_array[740] = 16'hbcbe;
mem_array[743] = 16'hd110;
mem_array[742] = 16'h3aca;
mem_array[745] = 16'hb716;
mem_array[744] = 16'hbd67;
mem_array[747] = 16'h5058;
mem_array[746] = 16'h3e27;
mem_array[749] = 16'h2f37;
mem_array[748] = 16'h3cfb;
mem_array[751] = 16'h304e;
mem_array[750] = 16'hbcef;
mem_array[753] = 16'he6e1;
mem_array[752] = 16'h3cba;
mem_array[755] = 16'hf540;
mem_array[754] = 16'hbd1b;
mem_array[757] = 16'hb86a;
mem_array[756] = 16'h3da7;
mem_array[759] = 16'hff55;
mem_array[758] = 16'hbd6b;
mem_array[761] = 16'h025a;
mem_array[760] = 16'h3d86;
mem_array[763] = 16'h10d5;
mem_array[762] = 16'hbdfe;
mem_array[765] = 16'h0afd;
mem_array[764] = 16'h3cc0;
mem_array[767] = 16'h0316;
mem_array[766] = 16'hbe1a;
mem_array[769] = 16'haec0;
mem_array[768] = 16'h3d7e;
mem_array[771] = 16'h14d9;
mem_array[770] = 16'h3cbb;
mem_array[773] = 16'h11ce;
mem_array[772] = 16'h3e1b;
mem_array[775] = 16'h0fa8;
mem_array[774] = 16'h3ccc;
mem_array[777] = 16'h8c60;
mem_array[776] = 16'h3b41;
mem_array[779] = 16'h9ea8;
mem_array[778] = 16'hbd8b;
mem_array[781] = 16'hd916;
mem_array[780] = 16'h3db2;
mem_array[783] = 16'h25ed;
mem_array[782] = 16'hbd3b;
mem_array[785] = 16'hc815;
mem_array[784] = 16'h3ca7;
mem_array[787] = 16'hefde;
mem_array[786] = 16'h3c6d;
mem_array[789] = 16'h2315;
mem_array[788] = 16'hbda9;
mem_array[791] = 16'h6f6b;
mem_array[790] = 16'h3c70;
mem_array[793] = 16'hc094;
mem_array[792] = 16'h3d86;
mem_array[795] = 16'hf35c;
mem_array[794] = 16'h3a0e;
mem_array[797] = 16'ha13a;
mem_array[796] = 16'h3d6a;
mem_array[799] = 16'he053;
mem_array[798] = 16'hbd43;
mem_array[801] = 16'hbe84;
mem_array[800] = 16'hbc03;
mem_array[803] = 16'ha4a3;
mem_array[802] = 16'h3db6;
mem_array[805] = 16'h85fe;
mem_array[804] = 16'h3bba;
mem_array[807] = 16'ha419;
mem_array[806] = 16'h3dfa;
mem_array[809] = 16'h8ea5;
mem_array[808] = 16'h3e1a;
mem_array[811] = 16'hfbc8;
mem_array[810] = 16'hbe51;
mem_array[813] = 16'h5cd9;
mem_array[812] = 16'hbd61;
mem_array[815] = 16'h0650;
mem_array[814] = 16'h3c75;
mem_array[817] = 16'h2c20;
mem_array[816] = 16'h3cdb;
mem_array[819] = 16'h540c;
mem_array[818] = 16'h3ceb;
mem_array[821] = 16'hd5ae;
mem_array[820] = 16'h3ca8;
mem_array[823] = 16'h1810;
mem_array[822] = 16'hbe29;
mem_array[825] = 16'hae13;
mem_array[824] = 16'h3d2d;
mem_array[827] = 16'h6aca;
mem_array[826] = 16'hbe85;
mem_array[829] = 16'hcd9b;
mem_array[828] = 16'h3e68;
mem_array[831] = 16'hbce8;
mem_array[830] = 16'h3d04;
mem_array[833] = 16'h32c1;
mem_array[832] = 16'h3e3b;
mem_array[835] = 16'h43f6;
mem_array[834] = 16'hbda1;
mem_array[837] = 16'hb1ef;
mem_array[836] = 16'h3e3b;
mem_array[839] = 16'hef4a;
mem_array[838] = 16'hbdcd;
mem_array[841] = 16'h19ca;
mem_array[840] = 16'hbcd0;
mem_array[843] = 16'h382f;
mem_array[842] = 16'hbcd6;
mem_array[845] = 16'he363;
mem_array[844] = 16'hbc11;
mem_array[847] = 16'h9ba6;
mem_array[846] = 16'h3c04;
mem_array[849] = 16'h0c1e;
mem_array[848] = 16'hbdb0;
mem_array[851] = 16'h8880;
mem_array[850] = 16'h3cfc;
mem_array[853] = 16'h1f76;
mem_array[852] = 16'hbd83;
mem_array[855] = 16'hf79e;
mem_array[854] = 16'h3d38;
mem_array[857] = 16'ha882;
mem_array[856] = 16'h3e21;
mem_array[859] = 16'hbb18;
mem_array[858] = 16'h3d4b;
mem_array[861] = 16'h3879;
mem_array[860] = 16'h3d22;
mem_array[863] = 16'h3f23;
mem_array[862] = 16'h3de1;
mem_array[865] = 16'hcc62;
mem_array[864] = 16'h39d5;
mem_array[867] = 16'h3fce;
mem_array[866] = 16'h3e15;
mem_array[869] = 16'h21b6;
mem_array[868] = 16'h3e66;
mem_array[871] = 16'h7444;
mem_array[870] = 16'hbe14;
mem_array[873] = 16'h9078;
mem_array[872] = 16'h3c95;
mem_array[875] = 16'h4d43;
mem_array[874] = 16'hbd55;
mem_array[877] = 16'h8d1e;
mem_array[876] = 16'hbd28;
mem_array[879] = 16'h44eb;
mem_array[878] = 16'hbc6d;
mem_array[881] = 16'h874b;
mem_array[880] = 16'hbdcb;
mem_array[883] = 16'hd1c5;
mem_array[882] = 16'hbe1e;
mem_array[885] = 16'h6626;
mem_array[884] = 16'hbd92;
mem_array[887] = 16'hfb2a;
mem_array[886] = 16'hbe6c;
mem_array[889] = 16'h2403;
mem_array[888] = 16'h3e5d;
mem_array[891] = 16'h4840;
mem_array[890] = 16'hbdb0;
mem_array[893] = 16'hca15;
mem_array[892] = 16'h3e33;
mem_array[895] = 16'he0d4;
mem_array[894] = 16'hbd0b;
mem_array[897] = 16'he0a2;
mem_array[896] = 16'h3ce0;
mem_array[899] = 16'h4540;
mem_array[898] = 16'hbc91;
mem_array[901] = 16'h0dad;
mem_array[900] = 16'h3d53;
mem_array[903] = 16'he32c;
mem_array[902] = 16'hbda1;
mem_array[905] = 16'hba56;
mem_array[904] = 16'hbc11;
mem_array[907] = 16'h6cf6;
mem_array[906] = 16'h3cda;
mem_array[909] = 16'he169;
mem_array[908] = 16'h3d00;
mem_array[911] = 16'h1f4f;
mem_array[910] = 16'h3d09;
mem_array[913] = 16'hc82e;
mem_array[912] = 16'hbd82;
mem_array[915] = 16'h4804;
mem_array[914] = 16'h3d2f;
mem_array[917] = 16'hd0f4;
mem_array[916] = 16'h3dea;
mem_array[919] = 16'hffbb;
mem_array[918] = 16'hbd5a;
mem_array[921] = 16'hf8b4;
mem_array[920] = 16'hbc8e;
mem_array[923] = 16'h212c;
mem_array[922] = 16'h3d7b;
mem_array[925] = 16'h5ba8;
mem_array[924] = 16'hbcbe;
mem_array[927] = 16'h6e04;
mem_array[926] = 16'h3de7;
mem_array[929] = 16'h8896;
mem_array[928] = 16'h3c28;
mem_array[931] = 16'he055;
mem_array[930] = 16'hbd55;
mem_array[933] = 16'hf44e;
mem_array[932] = 16'h3d7a;
mem_array[935] = 16'h5ac5;
mem_array[934] = 16'h3c87;
mem_array[937] = 16'h8a52;
mem_array[936] = 16'h3d9e;
mem_array[939] = 16'hc319;
mem_array[938] = 16'h3de0;
mem_array[941] = 16'h0055;
mem_array[940] = 16'hbcc3;
mem_array[943] = 16'hdb04;
mem_array[942] = 16'hbda7;
mem_array[945] = 16'h5f24;
mem_array[944] = 16'h3d84;
mem_array[947] = 16'hce63;
mem_array[946] = 16'hbe2b;
mem_array[949] = 16'h1e70;
mem_array[948] = 16'h3b82;
mem_array[951] = 16'h27e9;
mem_array[950] = 16'h3cba;
mem_array[953] = 16'h802d;
mem_array[952] = 16'h3d68;
mem_array[955] = 16'h27cf;
mem_array[954] = 16'h3d9c;
mem_array[957] = 16'h1897;
mem_array[956] = 16'h3bd9;
mem_array[959] = 16'ha49e;
mem_array[958] = 16'hbd20;
mem_array[961] = 16'h66eb;
mem_array[960] = 16'h3c79;
mem_array[963] = 16'hac45;
mem_array[962] = 16'hbd45;
mem_array[965] = 16'haaf3;
mem_array[964] = 16'hbd97;
mem_array[967] = 16'h106b;
mem_array[966] = 16'hbdce;
mem_array[969] = 16'h7e57;
mem_array[968] = 16'h3c82;
mem_array[971] = 16'h8324;
mem_array[970] = 16'hbd96;
mem_array[973] = 16'h2137;
mem_array[972] = 16'h3c55;
mem_array[975] = 16'h7959;
mem_array[974] = 16'h3d72;
mem_array[977] = 16'h4383;
mem_array[976] = 16'h3c3f;
mem_array[979] = 16'hc57f;
mem_array[978] = 16'hbd96;
mem_array[981] = 16'heffe;
mem_array[980] = 16'hbcec;
mem_array[983] = 16'h852e;
mem_array[982] = 16'h3db7;
mem_array[985] = 16'h84df;
mem_array[984] = 16'hbc9e;
mem_array[987] = 16'ha38c;
mem_array[986] = 16'h3dcd;
mem_array[989] = 16'h0b35;
mem_array[988] = 16'h3d46;
mem_array[991] = 16'h867f;
mem_array[990] = 16'h3d9c;
mem_array[993] = 16'h16bc;
mem_array[992] = 16'h3dde;
mem_array[995] = 16'h4055;
mem_array[994] = 16'h3c6a;
mem_array[997] = 16'h425c;
mem_array[996] = 16'h3d59;
mem_array[999] = 16'hfedd;
mem_array[998] = 16'h3d32;
mem_array[1001] = 16'h3ec0;
mem_array[1000] = 16'h3ce6;
mem_array[1003] = 16'h3239;
mem_array[1002] = 16'h3d01;
mem_array[1005] = 16'hfda4;
mem_array[1004] = 16'h3d6d;
mem_array[1007] = 16'h8cec;
mem_array[1006] = 16'h3d13;
mem_array[1009] = 16'h30e9;
mem_array[1008] = 16'h3cfb;
mem_array[1011] = 16'ha3dd;
mem_array[1010] = 16'hbd89;
mem_array[1013] = 16'hfeaf;
mem_array[1012] = 16'h3bfa;
mem_array[1015] = 16'hdde3;
mem_array[1014] = 16'h3d6d;
mem_array[1017] = 16'hf923;
mem_array[1016] = 16'hbcd5;
mem_array[1019] = 16'hdbdd;
mem_array[1018] = 16'hbc83;
mem_array[1021] = 16'hedae;
mem_array[1020] = 16'h3cde;
mem_array[1023] = 16'h4fb5;
mem_array[1022] = 16'hbd8b;
mem_array[1025] = 16'h5c99;
mem_array[1024] = 16'hbca6;
mem_array[1027] = 16'h36cb;
mem_array[1026] = 16'h3c69;
mem_array[1029] = 16'he99d;
mem_array[1028] = 16'hbbfc;
mem_array[1031] = 16'h3de1;
mem_array[1030] = 16'h3c7b;
mem_array[1033] = 16'h92b2;
mem_array[1032] = 16'hbd55;
mem_array[1035] = 16'hda4c;
mem_array[1034] = 16'hbbbb;
mem_array[1037] = 16'hcb4e;
mem_array[1036] = 16'hbcbb;
mem_array[1039] = 16'hed9b;
mem_array[1038] = 16'h3cc9;
mem_array[1041] = 16'hb3c7;
mem_array[1040] = 16'hbc14;
mem_array[1043] = 16'h1e96;
mem_array[1042] = 16'h3cdb;
mem_array[1045] = 16'h7159;
mem_array[1044] = 16'hbbae;
mem_array[1047] = 16'h107f;
mem_array[1046] = 16'h3d43;
mem_array[1049] = 16'hb3e4;
mem_array[1048] = 16'h3de8;
mem_array[1051] = 16'h0e96;
mem_array[1050] = 16'h3c0c;
mem_array[1053] = 16'heaf5;
mem_array[1052] = 16'h3caf;
mem_array[1055] = 16'h1566;
mem_array[1054] = 16'hbdbd;
mem_array[1057] = 16'h42b4;
mem_array[1056] = 16'h3b23;
mem_array[1059] = 16'hb34a;
mem_array[1058] = 16'hbdbe;
mem_array[1061] = 16'he92d;
mem_array[1060] = 16'hbd62;
mem_array[1063] = 16'h1658;
mem_array[1062] = 16'hbcaf;
mem_array[1065] = 16'he371;
mem_array[1064] = 16'hbcb8;
mem_array[1067] = 16'hece5;
mem_array[1066] = 16'hbd1f;
mem_array[1069] = 16'h75b1;
mem_array[1068] = 16'hbd3b;
mem_array[1071] = 16'h04c7;
mem_array[1070] = 16'h3cfa;
mem_array[1073] = 16'h6310;
mem_array[1072] = 16'hbd15;
mem_array[1075] = 16'ha790;
mem_array[1074] = 16'hbcbd;
mem_array[1077] = 16'he8d6;
mem_array[1076] = 16'hbd26;
mem_array[1079] = 16'h0c73;
mem_array[1078] = 16'hbcbe;
mem_array[1081] = 16'h516a;
mem_array[1080] = 16'hbcfa;
mem_array[1083] = 16'h0db2;
mem_array[1082] = 16'hbca4;
mem_array[1085] = 16'hf040;
mem_array[1084] = 16'hbcc5;
mem_array[1087] = 16'hfeb2;
mem_array[1086] = 16'h3d4e;
mem_array[1089] = 16'h9742;
mem_array[1088] = 16'hbcf4;
mem_array[1091] = 16'hc376;
mem_array[1090] = 16'h3b15;
mem_array[1093] = 16'hef06;
mem_array[1092] = 16'hbd8d;
mem_array[1095] = 16'hb94f;
mem_array[1094] = 16'h3c3f;
mem_array[1097] = 16'h3125;
mem_array[1096] = 16'hbd8d;
mem_array[1099] = 16'hea65;
mem_array[1098] = 16'hbb5a;
mem_array[1101] = 16'h1452;
mem_array[1100] = 16'h3d5f;
mem_array[1103] = 16'h64e5;
mem_array[1102] = 16'hbdbb;
mem_array[1105] = 16'hedcf;
mem_array[1104] = 16'hbd30;
mem_array[1107] = 16'h748f;
mem_array[1106] = 16'hbd62;
mem_array[1109] = 16'h8525;
mem_array[1108] = 16'h3d36;
mem_array[1111] = 16'hbfa2;
mem_array[1110] = 16'h3d00;
mem_array[1113] = 16'h6ad2;
mem_array[1112] = 16'h3d5f;
mem_array[1115] = 16'ha076;
mem_array[1114] = 16'hbc27;
mem_array[1117] = 16'h39d1;
mem_array[1116] = 16'h3d8e;
mem_array[1119] = 16'h9873;
mem_array[1118] = 16'hbc5b;
mem_array[1121] = 16'h0d36;
mem_array[1120] = 16'h3cb6;
mem_array[1123] = 16'h16ad;
mem_array[1122] = 16'hbdc0;
mem_array[1125] = 16'hf6d0;
mem_array[1124] = 16'hbb86;
mem_array[1127] = 16'h72d2;
mem_array[1126] = 16'hbd04;
mem_array[1129] = 16'hc924;
mem_array[1128] = 16'h3c19;
mem_array[1131] = 16'h7af8;
mem_array[1130] = 16'hbd49;
mem_array[1133] = 16'h34aa;
mem_array[1132] = 16'hbd4e;
mem_array[1135] = 16'hb6cf;
mem_array[1134] = 16'hbd71;
mem_array[1137] = 16'hadd8;
mem_array[1136] = 16'hbb6c;
mem_array[1139] = 16'h3baa;
mem_array[1138] = 16'hbc50;
mem_array[1141] = 16'hd34a;
mem_array[1140] = 16'h3bd4;
mem_array[1143] = 16'hf1c1;
mem_array[1142] = 16'hbb25;
mem_array[1145] = 16'h0b04;
mem_array[1144] = 16'h3c26;
mem_array[1147] = 16'h26dc;
mem_array[1146] = 16'h3d9a;
mem_array[1149] = 16'h6684;
mem_array[1148] = 16'h3c8a;
mem_array[1151] = 16'hd099;
mem_array[1150] = 16'hbd86;
mem_array[1153] = 16'h153e;
mem_array[1152] = 16'hbd99;
mem_array[1155] = 16'h5daf;
mem_array[1154] = 16'hbd56;
mem_array[1157] = 16'h1f81;
mem_array[1156] = 16'hbd67;
mem_array[1159] = 16'h7e45;
mem_array[1158] = 16'h3d64;
mem_array[1161] = 16'hafcf;
mem_array[1160] = 16'hbd44;
mem_array[1163] = 16'hd7f6;
mem_array[1162] = 16'hbd11;
mem_array[1165] = 16'h1759;
mem_array[1164] = 16'hbb27;
mem_array[1167] = 16'h7920;
mem_array[1166] = 16'hbd91;
mem_array[1169] = 16'hc2ec;
mem_array[1168] = 16'hbc9b;
mem_array[1171] = 16'hd64f;
mem_array[1170] = 16'hbbfd;
mem_array[1173] = 16'h2831;
mem_array[1172] = 16'h3c8f;
mem_array[1175] = 16'h300d;
mem_array[1174] = 16'h3dba;
mem_array[1177] = 16'h49ca;
mem_array[1176] = 16'h3d9d;
mem_array[1179] = 16'h6700;
mem_array[1178] = 16'h3d66;
mem_array[1181] = 16'h2948;
mem_array[1180] = 16'hbd25;
mem_array[1183] = 16'hc1fe;
mem_array[1182] = 16'hbdac;
mem_array[1185] = 16'h3ca7;
mem_array[1184] = 16'h3d32;
mem_array[1187] = 16'hb38e;
mem_array[1186] = 16'hbbb9;
mem_array[1189] = 16'h649a;
mem_array[1188] = 16'hbd27;
mem_array[1191] = 16'h757b;
mem_array[1190] = 16'h3d8f;
mem_array[1193] = 16'he2d0;
mem_array[1192] = 16'hbd46;
mem_array[1195] = 16'h2adf;
mem_array[1194] = 16'h3dad;
mem_array[1197] = 16'h0142;
mem_array[1196] = 16'hbd1a;
mem_array[1199] = 16'hd6da;
mem_array[1198] = 16'hbdb4;
mem_array[1201] = 16'h5267;
mem_array[1200] = 16'h3d11;
mem_array[1203] = 16'hc81d;
mem_array[1202] = 16'h3c65;
mem_array[1205] = 16'hab5f;
mem_array[1204] = 16'h3c8c;
mem_array[1207] = 16'hf9af;
mem_array[1206] = 16'hbd4f;
mem_array[1209] = 16'h21c9;
mem_array[1208] = 16'h3dcc;
mem_array[1211] = 16'h0190;
mem_array[1210] = 16'h3b5c;
mem_array[1213] = 16'ha54a;
mem_array[1212] = 16'hbd21;
mem_array[1215] = 16'h224a;
mem_array[1214] = 16'h3d4f;
mem_array[1217] = 16'h3ee2;
mem_array[1216] = 16'hbd01;
mem_array[1219] = 16'h853f;
mem_array[1218] = 16'hbcda;
mem_array[1221] = 16'hd42b;
mem_array[1220] = 16'hbd21;
mem_array[1223] = 16'h5720;
mem_array[1222] = 16'hba48;
mem_array[1225] = 16'h5682;
mem_array[1224] = 16'hbdd9;
mem_array[1227] = 16'h907b;
mem_array[1226] = 16'h3d32;
mem_array[1229] = 16'h4f67;
mem_array[1228] = 16'hbd98;
mem_array[1231] = 16'hfd62;
mem_array[1230] = 16'h3cea;
mem_array[1233] = 16'hc67b;
mem_array[1232] = 16'hbc9f;
mem_array[1235] = 16'h94f1;
mem_array[1234] = 16'h3be2;
mem_array[1237] = 16'h8a38;
mem_array[1236] = 16'h3d26;
mem_array[1239] = 16'h280a;
mem_array[1238] = 16'hbd78;
mem_array[1241] = 16'hcc32;
mem_array[1240] = 16'h3d19;
mem_array[1243] = 16'hec95;
mem_array[1242] = 16'h3c4f;
mem_array[1245] = 16'h27bf;
mem_array[1244] = 16'h3d11;
mem_array[1247] = 16'h4d54;
mem_array[1246] = 16'hbd5e;
mem_array[1249] = 16'habc6;
mem_array[1248] = 16'hbdbc;
mem_array[1251] = 16'hbab8;
mem_array[1250] = 16'h3c4b;
mem_array[1253] = 16'h0031;
mem_array[1252] = 16'h3dce;
mem_array[1255] = 16'hf07e;
mem_array[1254] = 16'h3a85;
mem_array[1257] = 16'h4bcd;
mem_array[1256] = 16'hbc8d;
mem_array[1259] = 16'h1531;
mem_array[1258] = 16'h3d0a;
mem_array[1261] = 16'hb492;
mem_array[1260] = 16'hbb87;
mem_array[1263] = 16'hb0ad;
mem_array[1262] = 16'h3d96;
mem_array[1265] = 16'hb66f;
mem_array[1264] = 16'h3c64;
mem_array[1267] = 16'h52cb;
mem_array[1266] = 16'h3d4a;
mem_array[1269] = 16'h26a7;
mem_array[1268] = 16'h3caf;
mem_array[1271] = 16'h91d6;
mem_array[1270] = 16'hbdd8;
mem_array[1273] = 16'h777b;
mem_array[1272] = 16'hbccb;
mem_array[1275] = 16'h26f7;
mem_array[1274] = 16'h3cd8;
mem_array[1277] = 16'hdd54;
mem_array[1276] = 16'hbd85;
mem_array[1279] = 16'h0776;
mem_array[1278] = 16'h3dc3;
mem_array[1281] = 16'hcbb4;
mem_array[1280] = 16'hbd29;
mem_array[1283] = 16'hb6f7;
mem_array[1282] = 16'hbc80;
mem_array[1285] = 16'h16b1;
mem_array[1284] = 16'hbd98;
mem_array[1287] = 16'h303d;
mem_array[1286] = 16'h3d86;
mem_array[1289] = 16'hcafc;
mem_array[1288] = 16'hbd31;
mem_array[1291] = 16'h8313;
mem_array[1290] = 16'h3c0f;
mem_array[1293] = 16'h6e8f;
mem_array[1292] = 16'h3bf5;
mem_array[1295] = 16'h6a68;
mem_array[1294] = 16'h3ceb;
mem_array[1297] = 16'heb65;
mem_array[1296] = 16'h3c54;
mem_array[1299] = 16'hb9b3;
mem_array[1298] = 16'h3d69;
mem_array[1301] = 16'h3108;
mem_array[1300] = 16'h3d64;
mem_array[1303] = 16'hb55f;
mem_array[1302] = 16'h3ce5;
mem_array[1305] = 16'h51de;
mem_array[1304] = 16'h3d4e;
mem_array[1307] = 16'ha9f5;
mem_array[1306] = 16'hbcbd;
mem_array[1309] = 16'hd4bc;
mem_array[1308] = 16'hbcb4;
mem_array[1311] = 16'ha178;
mem_array[1310] = 16'h3c4d;
mem_array[1313] = 16'hb7c2;
mem_array[1312] = 16'hbd0f;
mem_array[1315] = 16'h0705;
mem_array[1314] = 16'h3d4d;
mem_array[1317] = 16'h9243;
mem_array[1316] = 16'hbd69;
mem_array[1319] = 16'h2869;
mem_array[1318] = 16'h3d0d;
mem_array[1321] = 16'h4717;
mem_array[1320] = 16'hbd34;
mem_array[1323] = 16'h6eec;
mem_array[1322] = 16'hbcea;
mem_array[1325] = 16'h574c;
mem_array[1324] = 16'h3bdb;
mem_array[1327] = 16'h863d;
mem_array[1326] = 16'hbc64;
mem_array[1329] = 16'h55b7;
mem_array[1328] = 16'hbb4c;
mem_array[1331] = 16'h6873;
mem_array[1330] = 16'hbcab;
mem_array[1333] = 16'h883f;
mem_array[1332] = 16'h3cb0;
mem_array[1335] = 16'ha28f;
mem_array[1334] = 16'h3c00;
mem_array[1337] = 16'h8dcc;
mem_array[1336] = 16'h3cff;
mem_array[1339] = 16'h7878;
mem_array[1338] = 16'hbbeb;
mem_array[1341] = 16'h1746;
mem_array[1340] = 16'h3cb5;
mem_array[1343] = 16'h4070;
mem_array[1342] = 16'hbccd;
mem_array[1345] = 16'h6853;
mem_array[1344] = 16'hbd7a;
mem_array[1347] = 16'h1aea;
mem_array[1346] = 16'hbdd3;
mem_array[1349] = 16'h770d;
mem_array[1348] = 16'hbbef;
mem_array[1351] = 16'h8b51;
mem_array[1350] = 16'h3d4d;
mem_array[1353] = 16'h7472;
mem_array[1352] = 16'h3b8c;
mem_array[1355] = 16'h1c6e;
mem_array[1354] = 16'hbdc0;
mem_array[1357] = 16'he64c;
mem_array[1356] = 16'hbd36;
mem_array[1359] = 16'h88a7;
mem_array[1358] = 16'h3d22;
mem_array[1361] = 16'h3345;
mem_array[1360] = 16'h3d35;
mem_array[1363] = 16'h0d7d;
mem_array[1362] = 16'h3dc4;
mem_array[1365] = 16'h918e;
mem_array[1364] = 16'h3c24;
mem_array[1367] = 16'ha5b4;
mem_array[1366] = 16'hbd4b;
mem_array[1369] = 16'h09b7;
mem_array[1368] = 16'h3dde;
mem_array[1371] = 16'hc926;
mem_array[1370] = 16'hbc5b;
mem_array[1373] = 16'he371;
mem_array[1372] = 16'hbceb;
mem_array[1375] = 16'h1b81;
mem_array[1374] = 16'hbc86;
mem_array[1377] = 16'h23df;
mem_array[1376] = 16'hbd99;
mem_array[1379] = 16'h2619;
mem_array[1378] = 16'h3d9e;
mem_array[1381] = 16'h8fce;
mem_array[1380] = 16'hbc8e;
mem_array[1383] = 16'h0e6d;
mem_array[1382] = 16'h3a6c;
mem_array[1385] = 16'h3a58;
mem_array[1384] = 16'h3d26;
mem_array[1387] = 16'h3cff;
mem_array[1386] = 16'hbad0;
mem_array[1389] = 16'h8f49;
mem_array[1388] = 16'h3c88;
mem_array[1391] = 16'hbbbb;
mem_array[1390] = 16'hbd02;
mem_array[1393] = 16'h8e24;
mem_array[1392] = 16'hbd6f;
mem_array[1395] = 16'ha317;
mem_array[1394] = 16'hbd3b;
mem_array[1397] = 16'h70ad;
mem_array[1396] = 16'h3d91;
mem_array[1399] = 16'h2db7;
mem_array[1398] = 16'h3c96;
mem_array[1401] = 16'h12df;
mem_array[1400] = 16'hba94;
mem_array[1403] = 16'h80a7;
mem_array[1402] = 16'h3c8b;
mem_array[1405] = 16'hfaba;
mem_array[1404] = 16'h3c85;
mem_array[1407] = 16'hc6cc;
mem_array[1406] = 16'h3d7b;
mem_array[1409] = 16'ha3e1;
mem_array[1408] = 16'hbd25;
mem_array[1411] = 16'h3f06;
mem_array[1410] = 16'h3d20;
mem_array[1413] = 16'h92a9;
mem_array[1412] = 16'hbbd4;
mem_array[1415] = 16'hdeb9;
mem_array[1414] = 16'h3d7d;
mem_array[1417] = 16'h97d6;
mem_array[1416] = 16'h3da5;
mem_array[1419] = 16'ha7cb;
mem_array[1418] = 16'h3d3c;
mem_array[1421] = 16'h35e9;
mem_array[1420] = 16'hbda5;
mem_array[1423] = 16'h9dee;
mem_array[1422] = 16'h3d3f;
mem_array[1425] = 16'h42eb;
mem_array[1424] = 16'hbcb1;
mem_array[1427] = 16'h1533;
mem_array[1426] = 16'h3dc2;
mem_array[1429] = 16'h4f7d;
mem_array[1428] = 16'h3d11;
mem_array[1431] = 16'h1384;
mem_array[1430] = 16'hbd05;
mem_array[1433] = 16'h3a89;
mem_array[1432] = 16'h3cae;
mem_array[1435] = 16'h2b91;
mem_array[1434] = 16'h3d7f;
mem_array[1437] = 16'h449f;
mem_array[1436] = 16'hbca5;
mem_array[1439] = 16'hce81;
mem_array[1438] = 16'h3caf;
mem_array[1441] = 16'h1d4e;
mem_array[1440] = 16'hbcf2;
mem_array[1443] = 16'h28bd;
mem_array[1442] = 16'h3dcc;
mem_array[1445] = 16'hbfa6;
mem_array[1444] = 16'h3db6;
mem_array[1447] = 16'h349c;
mem_array[1446] = 16'h3bf4;
mem_array[1449] = 16'h2ad6;
mem_array[1448] = 16'h3d00;
mem_array[1451] = 16'hb306;
mem_array[1450] = 16'hbc5d;
mem_array[1453] = 16'hd63f;
mem_array[1452] = 16'hbab3;
mem_array[1455] = 16'h9b55;
mem_array[1454] = 16'hbc69;
mem_array[1457] = 16'h7eaf;
mem_array[1456] = 16'h3d23;
mem_array[1459] = 16'hca42;
mem_array[1458] = 16'hbcf2;
mem_array[1461] = 16'h420d;
mem_array[1460] = 16'h3d46;
mem_array[1463] = 16'h8a30;
mem_array[1462] = 16'hbd66;
mem_array[1465] = 16'hf62a;
mem_array[1464] = 16'hbd1f;
mem_array[1467] = 16'h0d0e;
mem_array[1466] = 16'hbb6f;
mem_array[1469] = 16'h561c;
mem_array[1468] = 16'h3d39;
mem_array[1471] = 16'h0854;
mem_array[1470] = 16'hbd17;
mem_array[1473] = 16'h0703;
mem_array[1472] = 16'hbd50;
mem_array[1475] = 16'h6bec;
mem_array[1474] = 16'h3dcd;
mem_array[1477] = 16'hfdba;
mem_array[1476] = 16'h3c7d;
mem_array[1479] = 16'hffc7;
mem_array[1478] = 16'hbcb6;
mem_array[1481] = 16'hd51b;
mem_array[1480] = 16'hbc34;
mem_array[1483] = 16'h25e4;
mem_array[1482] = 16'hbc00;
mem_array[1485] = 16'h4719;
mem_array[1484] = 16'hbc54;
mem_array[1487] = 16'h3686;
mem_array[1486] = 16'hbd9b;
mem_array[1489] = 16'h10e8;
mem_array[1488] = 16'h3c9d;
mem_array[1491] = 16'h9569;
mem_array[1490] = 16'h3abd;
mem_array[1493] = 16'hfd0e;
mem_array[1492] = 16'hbc05;
mem_array[1495] = 16'h3aef;
mem_array[1494] = 16'hbc94;
mem_array[1497] = 16'h9a7c;
mem_array[1496] = 16'h3c31;
mem_array[1499] = 16'h560e;
mem_array[1498] = 16'h3ccb;
mem_array[1501] = 16'h14d8;
mem_array[1500] = 16'h3ca0;
mem_array[1503] = 16'ha7f1;
mem_array[1502] = 16'h3d81;
mem_array[1505] = 16'h04bc;
mem_array[1504] = 16'h3c1b;
mem_array[1507] = 16'hc8a4;
mem_array[1506] = 16'hbc6b;
mem_array[1509] = 16'h566f;
mem_array[1508] = 16'hbd23;
mem_array[1511] = 16'h6dea;
mem_array[1510] = 16'hbdd2;
mem_array[1513] = 16'h940b;
mem_array[1512] = 16'hbc0f;
mem_array[1515] = 16'h5925;
mem_array[1514] = 16'hbc77;
mem_array[1517] = 16'h9615;
mem_array[1516] = 16'h3da9;
mem_array[1519] = 16'h74f7;
mem_array[1518] = 16'hbd31;
mem_array[1521] = 16'ha584;
mem_array[1520] = 16'h3d75;
mem_array[1523] = 16'h926c;
mem_array[1522] = 16'hbd86;
mem_array[1525] = 16'ha14d;
mem_array[1524] = 16'h3c7f;
mem_array[1527] = 16'h6b3f;
mem_array[1526] = 16'hbd18;
mem_array[1529] = 16'h0ed0;
mem_array[1528] = 16'h3d1d;
mem_array[1531] = 16'h4619;
mem_array[1530] = 16'h3d0b;
mem_array[1533] = 16'he89e;
mem_array[1532] = 16'h3d20;
mem_array[1535] = 16'h4897;
mem_array[1534] = 16'hbd99;
mem_array[1537] = 16'h8456;
mem_array[1536] = 16'hbc71;
mem_array[1539] = 16'hca03;
mem_array[1538] = 16'h3c34;
mem_array[1541] = 16'h8697;
mem_array[1540] = 16'h3cc6;
mem_array[1543] = 16'hf393;
mem_array[1542] = 16'hbd02;
mem_array[1545] = 16'h7a02;
mem_array[1544] = 16'hbca9;
mem_array[1547] = 16'h527a;
mem_array[1546] = 16'hbd9a;
mem_array[1549] = 16'h4d54;
mem_array[1548] = 16'h3d0f;
mem_array[1551] = 16'h03c5;
mem_array[1550] = 16'h3dd8;
mem_array[1553] = 16'h7719;
mem_array[1552] = 16'hbd94;
mem_array[1555] = 16'hfe16;
mem_array[1554] = 16'hbd52;
mem_array[1557] = 16'hdd5a;
mem_array[1556] = 16'hbdc9;
mem_array[1559] = 16'ha14b;
mem_array[1558] = 16'h3cb9;
mem_array[1561] = 16'hbc99;
mem_array[1560] = 16'h3daa;
mem_array[1563] = 16'he75a;
mem_array[1562] = 16'h3cd0;
mem_array[1565] = 16'h8d75;
mem_array[1564] = 16'hbc50;
mem_array[1567] = 16'h7def;
mem_array[1566] = 16'hbc27;
mem_array[1569] = 16'h7459;
mem_array[1568] = 16'h3bf4;
mem_array[1571] = 16'hce99;
mem_array[1570] = 16'hbb9f;
mem_array[1573] = 16'hddba;
mem_array[1572] = 16'hbd61;
mem_array[1575] = 16'hefac;
mem_array[1574] = 16'h3d2e;
mem_array[1577] = 16'hd627;
mem_array[1576] = 16'hbc18;
mem_array[1579] = 16'ha2dd;
mem_array[1578] = 16'h3c89;
mem_array[1581] = 16'hbc89;
mem_array[1580] = 16'h3cb1;
mem_array[1583] = 16'h828e;
mem_array[1582] = 16'h3cdf;
mem_array[1585] = 16'h5048;
mem_array[1584] = 16'h3d6a;
mem_array[1587] = 16'h5419;
mem_array[1586] = 16'h3d21;
mem_array[1589] = 16'hd48e;
mem_array[1588] = 16'h3da5;
mem_array[1591] = 16'h6f35;
mem_array[1590] = 16'hbc79;
mem_array[1593] = 16'h28bd;
mem_array[1592] = 16'h3dbd;
mem_array[1595] = 16'h04b8;
mem_array[1594] = 16'h3bd8;
mem_array[1597] = 16'h5df9;
mem_array[1596] = 16'hbb75;
mem_array[1599] = 16'ha12b;
mem_array[1598] = 16'h3d8c;
mem_array[1601] = 16'h4daa;
mem_array[1600] = 16'hba92;
mem_array[1603] = 16'hb249;
mem_array[1602] = 16'hbd22;
mem_array[1605] = 16'h94fd;
mem_array[1604] = 16'hbd75;
mem_array[1607] = 16'h4124;
mem_array[1606] = 16'hbc39;
mem_array[1609] = 16'hd32a;
mem_array[1608] = 16'hbd2e;
mem_array[1611] = 16'h0063;
mem_array[1610] = 16'h3d7f;
mem_array[1613] = 16'h0ad0;
mem_array[1612] = 16'hbd17;
mem_array[1615] = 16'hbdc2;
mem_array[1614] = 16'h3d77;
mem_array[1617] = 16'h259a;
mem_array[1616] = 16'hbdaf;
mem_array[1619] = 16'h9341;
mem_array[1618] = 16'hbdd9;
mem_array[1621] = 16'hb33f;
mem_array[1620] = 16'hbd23;
mem_array[1623] = 16'h20e1;
mem_array[1622] = 16'h3d3e;
mem_array[1625] = 16'h6ada;
mem_array[1624] = 16'hbd81;
mem_array[1627] = 16'h7f2c;
mem_array[1626] = 16'h3ab6;
mem_array[1629] = 16'h5df8;
mem_array[1628] = 16'h3d3f;
mem_array[1631] = 16'h9a1d;
mem_array[1630] = 16'h3c43;
mem_array[1633] = 16'h899d;
mem_array[1632] = 16'h3cbd;
mem_array[1635] = 16'h4b72;
mem_array[1634] = 16'hbcb0;
mem_array[1637] = 16'h2dd0;
mem_array[1636] = 16'hbcad;
mem_array[1639] = 16'hd60c;
mem_array[1638] = 16'hbd3f;
mem_array[1641] = 16'hf957;
mem_array[1640] = 16'hbd03;
mem_array[1643] = 16'h83c4;
mem_array[1642] = 16'h3d80;
mem_array[1645] = 16'h23bf;
mem_array[1644] = 16'hbd10;
mem_array[1647] = 16'hc925;
mem_array[1646] = 16'h3d93;
mem_array[1649] = 16'h077e;
mem_array[1648] = 16'h3d3f;
mem_array[1651] = 16'hb515;
mem_array[1650] = 16'hbcce;
mem_array[1653] = 16'h33f4;
mem_array[1652] = 16'hbdac;
mem_array[1655] = 16'hd20f;
mem_array[1654] = 16'hbd13;
mem_array[1657] = 16'he2f0;
mem_array[1656] = 16'hbc8e;
mem_array[1659] = 16'h3573;
mem_array[1658] = 16'hbca3;
mem_array[1661] = 16'hfa28;
mem_array[1660] = 16'hbdbe;
mem_array[1663] = 16'h67fc;
mem_array[1662] = 16'hbd72;
mem_array[1665] = 16'h1ffb;
mem_array[1664] = 16'hbd17;
mem_array[1667] = 16'h1c8a;
mem_array[1666] = 16'hbcd2;
mem_array[1669] = 16'hf0c3;
mem_array[1668] = 16'hbd57;
mem_array[1671] = 16'he136;
mem_array[1670] = 16'hbd54;
mem_array[1673] = 16'he526;
mem_array[1672] = 16'hbd44;
mem_array[1675] = 16'h18e6;
mem_array[1674] = 16'hbb74;
mem_array[1677] = 16'h9871;
mem_array[1676] = 16'hbddc;
mem_array[1679] = 16'hc8f1;
mem_array[1678] = 16'hbd07;
mem_array[1681] = 16'h7482;
mem_array[1680] = 16'h3d21;
mem_array[1683] = 16'hb472;
mem_array[1682] = 16'h3d5c;
mem_array[1685] = 16'hfb82;
mem_array[1684] = 16'hbc34;
mem_array[1687] = 16'h6051;
mem_array[1686] = 16'h3d51;
mem_array[1689] = 16'hc33b;
mem_array[1688] = 16'h3d61;
mem_array[1691] = 16'h4258;
mem_array[1690] = 16'h3dbe;
mem_array[1693] = 16'h33a8;
mem_array[1692] = 16'h3d85;
mem_array[1695] = 16'h37fb;
mem_array[1694] = 16'hbdb2;
mem_array[1697] = 16'h7ddc;
mem_array[1696] = 16'hb963;
mem_array[1699] = 16'h39a0;
mem_array[1698] = 16'hbd72;
mem_array[1701] = 16'h74d3;
mem_array[1700] = 16'h3d61;
mem_array[1703] = 16'hcd6d;
mem_array[1702] = 16'h3d3b;
mem_array[1705] = 16'ha41d;
mem_array[1704] = 16'hbcbe;
mem_array[1707] = 16'hed8c;
mem_array[1706] = 16'hbd5f;
mem_array[1709] = 16'h4c5f;
mem_array[1708] = 16'hbd2b;
mem_array[1711] = 16'h6d57;
mem_array[1710] = 16'hbcf7;
mem_array[1713] = 16'hcaec;
mem_array[1712] = 16'h3b33;
mem_array[1715] = 16'hb334;
mem_array[1714] = 16'h3c0c;
mem_array[1717] = 16'h5361;
mem_array[1716] = 16'h3d20;
mem_array[1719] = 16'hc5bb;
mem_array[1718] = 16'hbcbe;
mem_array[1721] = 16'h0a3c;
mem_array[1720] = 16'h3cb7;
mem_array[1723] = 16'h1e2b;
mem_array[1722] = 16'h3cdb;
mem_array[1725] = 16'h88d9;
mem_array[1724] = 16'h3ddb;
mem_array[1727] = 16'h091c;
mem_array[1726] = 16'h3d65;
mem_array[1729] = 16'h78e1;
mem_array[1728] = 16'h3dc4;
mem_array[1731] = 16'h382b;
mem_array[1730] = 16'h3d29;
mem_array[1733] = 16'h15fc;
mem_array[1732] = 16'hbd08;
mem_array[1735] = 16'h5bf8;
mem_array[1734] = 16'h3c6d;
mem_array[1737] = 16'h695d;
mem_array[1736] = 16'h3daf;
mem_array[1739] = 16'h5300;
mem_array[1738] = 16'hbc82;
mem_array[1741] = 16'hce29;
mem_array[1740] = 16'h3da4;
mem_array[1743] = 16'h1f3e;
mem_array[1742] = 16'hbcc7;
mem_array[1745] = 16'h41fb;
mem_array[1744] = 16'hbd23;
mem_array[1747] = 16'h0659;
mem_array[1746] = 16'h3994;
mem_array[1749] = 16'h05b5;
mem_array[1748] = 16'hbc7c;
mem_array[1751] = 16'hc42c;
mem_array[1750] = 16'hbc59;
mem_array[1753] = 16'h6b7f;
mem_array[1752] = 16'hbc1b;
mem_array[1755] = 16'h7476;
mem_array[1754] = 16'h3d87;
mem_array[1757] = 16'heb40;
mem_array[1756] = 16'h3db1;
mem_array[1759] = 16'h696d;
mem_array[1758] = 16'hbdb6;
mem_array[1761] = 16'hf87a;
mem_array[1760] = 16'h3d25;
mem_array[1763] = 16'h8bc7;
mem_array[1762] = 16'h3da6;
mem_array[1765] = 16'ha891;
mem_array[1764] = 16'h3d75;
mem_array[1767] = 16'he1d4;
mem_array[1766] = 16'h3cd8;
mem_array[1769] = 16'h1736;
mem_array[1768] = 16'h3d20;
mem_array[1771] = 16'h8b3a;
mem_array[1770] = 16'h3d21;
mem_array[1773] = 16'hc661;
mem_array[1772] = 16'hbcdb;
mem_array[1775] = 16'h0cc1;
mem_array[1774] = 16'hbdbf;
mem_array[1777] = 16'h1041;
mem_array[1776] = 16'hbcf8;
mem_array[1779] = 16'h059c;
mem_array[1778] = 16'hbd65;
mem_array[1781] = 16'h98bd;
mem_array[1780] = 16'h3d19;
mem_array[1783] = 16'hf5f0;
mem_array[1782] = 16'h3d35;
mem_array[1785] = 16'haeca;
mem_array[1784] = 16'h3dc4;
mem_array[1787] = 16'h384b;
mem_array[1786] = 16'h3d11;
mem_array[1789] = 16'h7a0c;
mem_array[1788] = 16'hbd37;
mem_array[1791] = 16'h3e0c;
mem_array[1790] = 16'hbbcf;
mem_array[1793] = 16'hca83;
mem_array[1792] = 16'hbcbc;
mem_array[1795] = 16'h1625;
mem_array[1794] = 16'h3d40;
mem_array[1797] = 16'h4366;
mem_array[1796] = 16'hbd23;
mem_array[1799] = 16'h24de;
mem_array[1798] = 16'h3c8d;
mem_array[1801] = 16'h0145;
mem_array[1800] = 16'h3ca2;
mem_array[1803] = 16'h0ac3;
mem_array[1802] = 16'hbcae;
mem_array[1805] = 16'h85a4;
mem_array[1804] = 16'h3d30;
mem_array[1807] = 16'h6fc1;
mem_array[1806] = 16'hbca3;
mem_array[1809] = 16'h80b9;
mem_array[1808] = 16'hbd8a;
mem_array[1811] = 16'he0aa;
mem_array[1810] = 16'h3d98;
mem_array[1813] = 16'h5e83;
mem_array[1812] = 16'hbc8b;
mem_array[1815] = 16'h1fb3;
mem_array[1814] = 16'h3c0d;
mem_array[1817] = 16'ha05c;
mem_array[1816] = 16'hbb98;
mem_array[1819] = 16'hc03b;
mem_array[1818] = 16'h3c8f;
mem_array[1821] = 16'hf38a;
mem_array[1820] = 16'h3d23;
mem_array[1823] = 16'h99a8;
mem_array[1822] = 16'hbd23;
mem_array[1825] = 16'h7e56;
mem_array[1824] = 16'h3d31;
mem_array[1827] = 16'h6888;
mem_array[1826] = 16'hbcef;
mem_array[1829] = 16'h5fef;
mem_array[1828] = 16'h3c6a;
mem_array[1831] = 16'h3f25;
mem_array[1830] = 16'hbc31;
mem_array[1833] = 16'h059e;
mem_array[1832] = 16'hbcd9;
mem_array[1835] = 16'h6b90;
mem_array[1834] = 16'h3c67;
mem_array[1837] = 16'h58f7;
mem_array[1836] = 16'h3d3a;
mem_array[1839] = 16'h323a;
mem_array[1838] = 16'hbcb9;
mem_array[1841] = 16'h2add;
mem_array[1840] = 16'h3b3d;
mem_array[1843] = 16'h7c16;
mem_array[1842] = 16'hbdc7;
mem_array[1845] = 16'h128d;
mem_array[1844] = 16'hbcb2;
mem_array[1847] = 16'h0bb3;
mem_array[1846] = 16'h3a69;
mem_array[1849] = 16'h7396;
mem_array[1848] = 16'h3d16;
mem_array[1851] = 16'hb862;
mem_array[1850] = 16'h3cf3;
mem_array[1853] = 16'he147;
mem_array[1852] = 16'h3da3;
mem_array[1855] = 16'h38e8;
mem_array[1854] = 16'h3d30;
mem_array[1857] = 16'h4f61;
mem_array[1856] = 16'h3c1f;
mem_array[1859] = 16'h976b;
mem_array[1858] = 16'h3de7;
mem_array[1861] = 16'h94f0;
mem_array[1860] = 16'h3c88;
mem_array[1863] = 16'he470;
mem_array[1862] = 16'hbb60;
mem_array[1865] = 16'hf5f2;
mem_array[1864] = 16'h3dac;
mem_array[1867] = 16'he3c3;
mem_array[1866] = 16'h3cda;
mem_array[1869] = 16'h277f;
mem_array[1868] = 16'h3c88;
mem_array[1871] = 16'h006c;
mem_array[1870] = 16'h3d1c;
mem_array[1873] = 16'h8ae6;
mem_array[1872] = 16'hbdb6;
mem_array[1875] = 16'hd698;
mem_array[1874] = 16'h3d45;
mem_array[1877] = 16'he14e;
mem_array[1876] = 16'hbd50;
mem_array[1879] = 16'h3961;
mem_array[1878] = 16'hbd5c;
mem_array[1881] = 16'hf790;
mem_array[1880] = 16'hbb2f;
mem_array[1883] = 16'h3901;
mem_array[1882] = 16'h3d27;
mem_array[1885] = 16'h552f;
mem_array[1884] = 16'h3c73;
mem_array[1887] = 16'h7016;
mem_array[1886] = 16'hbde4;
mem_array[1889] = 16'h41a1;
mem_array[1888] = 16'hbd85;
mem_array[1891] = 16'h10c0;
mem_array[1890] = 16'hbd34;
mem_array[1893] = 16'h6340;
mem_array[1892] = 16'h3c8f;
mem_array[1895] = 16'h81b0;
mem_array[1894] = 16'h3dae;
mem_array[1897] = 16'h68a3;
mem_array[1896] = 16'h3c7d;
mem_array[1899] = 16'h29ea;
mem_array[1898] = 16'hbcac;
mem_array[1901] = 16'hf763;
mem_array[1900] = 16'hbcc0;
mem_array[1903] = 16'h97df;
mem_array[1902] = 16'h3c97;
mem_array[1905] = 16'heb50;
mem_array[1904] = 16'hbdcd;
mem_array[1907] = 16'hace7;
mem_array[1906] = 16'hbb88;
mem_array[1909] = 16'h533d;
mem_array[1908] = 16'h3c9a;
mem_array[1911] = 16'h98ba;
mem_array[1910] = 16'hbbcd;
mem_array[1913] = 16'h415d;
mem_array[1912] = 16'h3d77;
mem_array[1915] = 16'h8941;
mem_array[1914] = 16'h3d11;
mem_array[1917] = 16'hc952;
mem_array[1916] = 16'h3d45;
mem_array[1919] = 16'h3289;
mem_array[1918] = 16'h3dcb;
mem_array[1921] = 16'h8866;
mem_array[1920] = 16'hbd2a;
mem_array[1923] = 16'h69d7;
mem_array[1922] = 16'h3d48;
mem_array[1925] = 16'h168c;
mem_array[1924] = 16'hbdb3;
mem_array[1927] = 16'hea44;
mem_array[1926] = 16'h3c89;
mem_array[1929] = 16'h2e5b;
mem_array[1928] = 16'hbde4;
mem_array[1931] = 16'hd07d;
mem_array[1930] = 16'h3da6;
mem_array[1933] = 16'hb8e6;
mem_array[1932] = 16'hbd79;
mem_array[1935] = 16'hc891;
mem_array[1934] = 16'hbcc1;
mem_array[1937] = 16'h17c1;
mem_array[1936] = 16'hbcdc;
mem_array[1939] = 16'h9edf;
mem_array[1938] = 16'h3d53;
mem_array[1941] = 16'h399d;
mem_array[1940] = 16'hbbc2;
mem_array[1943] = 16'h12c2;
mem_array[1942] = 16'hbd35;
mem_array[1945] = 16'h5726;
mem_array[1944] = 16'h3cda;
mem_array[1947] = 16'h42a6;
mem_array[1946] = 16'h3c88;
mem_array[1949] = 16'h53df;
mem_array[1948] = 16'h3d2b;
mem_array[1951] = 16'h2613;
mem_array[1950] = 16'hbcda;
mem_array[1953] = 16'h6ab4;
mem_array[1952] = 16'hbb01;
mem_array[1955] = 16'h0ddd;
mem_array[1954] = 16'hbd8a;
mem_array[1957] = 16'he027;
mem_array[1956] = 16'hbcc7;
mem_array[1959] = 16'hdca9;
mem_array[1958] = 16'hbd07;
mem_array[1961] = 16'h9915;
mem_array[1960] = 16'hbc55;
mem_array[1963] = 16'hcb99;
mem_array[1962] = 16'h3d4b;
mem_array[1965] = 16'h8b06;
mem_array[1964] = 16'hbd26;
mem_array[1967] = 16'h5392;
mem_array[1966] = 16'h3d4c;
mem_array[1969] = 16'h3ddf;
mem_array[1968] = 16'h3ddd;
mem_array[1971] = 16'hd229;
mem_array[1970] = 16'h3ad7;
mem_array[1973] = 16'hafdd;
mem_array[1972] = 16'hbcfe;
mem_array[1975] = 16'h399a;
mem_array[1974] = 16'hbc06;
mem_array[1977] = 16'hac6e;
mem_array[1976] = 16'h3d40;
mem_array[1979] = 16'he2bb;
mem_array[1978] = 16'h3cd0;
mem_array[1981] = 16'h3210;
mem_array[1980] = 16'hbc85;
mem_array[1983] = 16'h3f76;
mem_array[1982] = 16'hbd98;
mem_array[1985] = 16'h6b40;
mem_array[1984] = 16'hbd49;
mem_array[1987] = 16'h2f0e;
mem_array[1986] = 16'h3d50;
mem_array[1989] = 16'haf6b;
mem_array[1988] = 16'h3d91;
mem_array[1991] = 16'h33ed;
mem_array[1990] = 16'h3d78;
mem_array[1993] = 16'h182a;
mem_array[1992] = 16'h3cd2;
mem_array[1995] = 16'h2ad2;
mem_array[1994] = 16'hbd55;
mem_array[1997] = 16'ha329;
mem_array[1996] = 16'hbc76;
mem_array[1999] = 16'hd04d;
mem_array[1998] = 16'h3c44;
mem_array[2001] = 16'hb9df;
mem_array[2000] = 16'h3cc7;
mem_array[2003] = 16'hc0b1;
mem_array[2002] = 16'h3d45;
mem_array[2005] = 16'hac0f;
mem_array[2004] = 16'h3def;
mem_array[2007] = 16'he13b;
mem_array[2006] = 16'h3c97;
mem_array[2009] = 16'hca1a;
mem_array[2008] = 16'hbdae;
mem_array[2011] = 16'h56ad;
mem_array[2010] = 16'hbdbe;
mem_array[2013] = 16'he1e7;
mem_array[2012] = 16'hbb64;
mem_array[2015] = 16'h7f32;
mem_array[2014] = 16'hbbb9;
mem_array[2017] = 16'hf37f;
mem_array[2016] = 16'h3cff;
mem_array[2019] = 16'h8a12;
mem_array[2018] = 16'hbd6d;
mem_array[2021] = 16'h490f;
mem_array[2020] = 16'h3d1d;
mem_array[2023] = 16'hf3b1;
mem_array[2022] = 16'h3dc3;
mem_array[2025] = 16'h39c6;
mem_array[2024] = 16'h3d01;
mem_array[2027] = 16'h4ff8;
mem_array[2026] = 16'h3d8f;
mem_array[2029] = 16'h273b;
mem_array[2028] = 16'hbde7;
mem_array[2031] = 16'hffc4;
mem_array[2030] = 16'h3b92;
mem_array[2033] = 16'h4f8e;
mem_array[2032] = 16'h3d80;
mem_array[2035] = 16'hfd95;
mem_array[2034] = 16'h3d76;
mem_array[2037] = 16'hfbf2;
mem_array[2036] = 16'hbd3e;
mem_array[2039] = 16'h8ae2;
mem_array[2038] = 16'hbdf2;
mem_array[2041] = 16'h9291;
mem_array[2040] = 16'hbd33;
mem_array[2043] = 16'h12b9;
mem_array[2042] = 16'hbb4a;
mem_array[2045] = 16'hae7d;
mem_array[2044] = 16'h3d4e;
mem_array[2047] = 16'ha4fa;
mem_array[2046] = 16'hbd50;
mem_array[2049] = 16'hbf60;
mem_array[2048] = 16'hbd13;
mem_array[2051] = 16'h30e5;
mem_array[2050] = 16'hbdd8;
mem_array[2053] = 16'h80d5;
mem_array[2052] = 16'hbe0a;
mem_array[2055] = 16'ha054;
mem_array[2054] = 16'h3d37;
mem_array[2057] = 16'h7117;
mem_array[2056] = 16'hbe80;
mem_array[2059] = 16'hac56;
mem_array[2058] = 16'h3c7d;
mem_array[2061] = 16'hf32c;
mem_array[2060] = 16'h3b7d;
mem_array[2063] = 16'h3eaf;
mem_array[2062] = 16'hbd4b;
mem_array[2065] = 16'h0308;
mem_array[2064] = 16'h3e69;
mem_array[2067] = 16'ha366;
mem_array[2066] = 16'hbc83;
mem_array[2069] = 16'hfd54;
mem_array[2068] = 16'hbd3f;
mem_array[2071] = 16'h9650;
mem_array[2070] = 16'h3d86;
mem_array[2073] = 16'hcf04;
mem_array[2072] = 16'hbd90;
mem_array[2075] = 16'hd068;
mem_array[2074] = 16'hbd80;
mem_array[2077] = 16'h18cb;
mem_array[2076] = 16'hbe63;
mem_array[2079] = 16'h32a2;
mem_array[2078] = 16'hbecb;
mem_array[2081] = 16'hacc7;
mem_array[2080] = 16'hbdc2;
mem_array[2083] = 16'h807e;
mem_array[2082] = 16'h3efc;
mem_array[2085] = 16'hadc5;
mem_array[2084] = 16'hbd95;
mem_array[2087] = 16'h6eaa;
mem_array[2086] = 16'h3ecb;
mem_array[2089] = 16'hc41f;
mem_array[2088] = 16'hbdc9;
mem_array[2091] = 16'h2c94;
mem_array[2090] = 16'hbe25;
mem_array[2093] = 16'ha464;
mem_array[2092] = 16'h3e6f;
mem_array[2095] = 16'h8a50;
mem_array[2094] = 16'h3d9a;
mem_array[2097] = 16'he856;
mem_array[2096] = 16'hbd9e;
mem_array[2099] = 16'hbef7;
mem_array[2098] = 16'hbe5e;
mem_array[2101] = 16'hce9c;
mem_array[2100] = 16'h3d89;
mem_array[2103] = 16'h3fb1;
mem_array[2102] = 16'h3c75;
mem_array[2105] = 16'h7740;
mem_array[2104] = 16'h3a37;
mem_array[2107] = 16'h8528;
mem_array[2106] = 16'hbcbb;
mem_array[2109] = 16'h8ce5;
mem_array[2108] = 16'hbd8b;
mem_array[2111] = 16'h14e3;
mem_array[2110] = 16'hbcb3;
mem_array[2113] = 16'h64a3;
mem_array[2112] = 16'hbd2d;
mem_array[2115] = 16'ha804;
mem_array[2114] = 16'h3cce;
mem_array[2117] = 16'hd45b;
mem_array[2116] = 16'hbea4;
mem_array[2119] = 16'hf7ef;
mem_array[2118] = 16'h3a02;
mem_array[2121] = 16'h5c86;
mem_array[2120] = 16'hbdcc;
mem_array[2123] = 16'hc337;
mem_array[2122] = 16'hbd72;
mem_array[2125] = 16'hc1c6;
mem_array[2124] = 16'h3e93;
mem_array[2127] = 16'h6c97;
mem_array[2126] = 16'hbc8c;
mem_array[2129] = 16'h6e16;
mem_array[2128] = 16'h3d43;
mem_array[2131] = 16'ha15c;
mem_array[2130] = 16'h3bb6;
mem_array[2133] = 16'h566f;
mem_array[2132] = 16'h3e00;
mem_array[2135] = 16'hd67e;
mem_array[2134] = 16'hbdf9;
mem_array[2137] = 16'ha517;
mem_array[2136] = 16'hbe8c;
mem_array[2139] = 16'h2903;
mem_array[2138] = 16'hbec5;
mem_array[2141] = 16'h7abd;
mem_array[2140] = 16'hbe1e;
mem_array[2143] = 16'hff9c;
mem_array[2142] = 16'h3ead;
mem_array[2145] = 16'ha476;
mem_array[2144] = 16'h3d5b;
mem_array[2147] = 16'h60f7;
mem_array[2146] = 16'h3ef8;
mem_array[2149] = 16'h7db6;
mem_array[2148] = 16'hbdad;
mem_array[2151] = 16'hfc55;
mem_array[2150] = 16'hbca7;
mem_array[2153] = 16'h6659;
mem_array[2152] = 16'h3c89;
mem_array[2155] = 16'hc077;
mem_array[2154] = 16'h3d0e;
mem_array[2157] = 16'hc042;
mem_array[2156] = 16'hbe78;
mem_array[2159] = 16'h2293;
mem_array[2158] = 16'hbe27;
mem_array[2161] = 16'hab17;
mem_array[2160] = 16'h3daf;
mem_array[2163] = 16'h9399;
mem_array[2162] = 16'hbd39;
mem_array[2165] = 16'h51ee;
mem_array[2164] = 16'hbd55;
mem_array[2167] = 16'hdda8;
mem_array[2166] = 16'h3e17;
mem_array[2169] = 16'hbdde;
mem_array[2168] = 16'hbea6;
mem_array[2171] = 16'h5739;
mem_array[2170] = 16'h3d71;
mem_array[2173] = 16'h7bf3;
mem_array[2172] = 16'hbee9;
mem_array[2175] = 16'h22a2;
mem_array[2174] = 16'h3dff;
mem_array[2177] = 16'h253a;
mem_array[2176] = 16'hbdf2;
mem_array[2179] = 16'h8ce8;
mem_array[2178] = 16'hba43;
mem_array[2181] = 16'h004d;
mem_array[2180] = 16'hbd15;
mem_array[2183] = 16'h0eb4;
mem_array[2182] = 16'hbcaf;
mem_array[2185] = 16'hf7a7;
mem_array[2184] = 16'h3f15;
mem_array[2187] = 16'h0490;
mem_array[2186] = 16'hbdee;
mem_array[2189] = 16'h6c85;
mem_array[2188] = 16'h3cb7;
mem_array[2191] = 16'hc901;
mem_array[2190] = 16'hbd8b;
mem_array[2193] = 16'h6304;
mem_array[2192] = 16'h3d8a;
mem_array[2195] = 16'h70cb;
mem_array[2194] = 16'hbdce;
mem_array[2197] = 16'hcbfc;
mem_array[2196] = 16'hbde2;
mem_array[2199] = 16'h8d92;
mem_array[2198] = 16'hbe7c;
mem_array[2201] = 16'h26da;
mem_array[2200] = 16'hbde4;
mem_array[2203] = 16'hb306;
mem_array[2202] = 16'hbc85;
mem_array[2205] = 16'h0d88;
mem_array[2204] = 16'hbe22;
mem_array[2207] = 16'ha1bb;
mem_array[2206] = 16'h3f35;
mem_array[2209] = 16'h3f8a;
mem_array[2208] = 16'hbdd0;
mem_array[2211] = 16'h24ff;
mem_array[2210] = 16'hbd03;
mem_array[2213] = 16'h27be;
mem_array[2212] = 16'hbe46;
mem_array[2215] = 16'hea3e;
mem_array[2214] = 16'h3ce2;
mem_array[2217] = 16'h242f;
mem_array[2216] = 16'hbdb0;
mem_array[2219] = 16'h3419;
mem_array[2218] = 16'hbdc6;
mem_array[2221] = 16'he1ed;
mem_array[2220] = 16'h3d0f;
mem_array[2223] = 16'h7c80;
mem_array[2222] = 16'hbd1e;
mem_array[2225] = 16'hd95b;
mem_array[2224] = 16'hbc6f;
mem_array[2227] = 16'h6ddb;
mem_array[2226] = 16'h3f5a;
mem_array[2229] = 16'h00dd;
mem_array[2228] = 16'hbef1;
mem_array[2231] = 16'h8a07;
mem_array[2230] = 16'h3d6d;
mem_array[2233] = 16'hb745;
mem_array[2232] = 16'hbfaa;
mem_array[2235] = 16'hea4b;
mem_array[2234] = 16'h3db3;
mem_array[2237] = 16'h5f3c;
mem_array[2236] = 16'hbeba;
mem_array[2239] = 16'h9543;
mem_array[2238] = 16'hbde1;
mem_array[2241] = 16'h83dc;
mem_array[2240] = 16'hbc8f;
mem_array[2243] = 16'h6438;
mem_array[2242] = 16'h3ccb;
mem_array[2245] = 16'hd807;
mem_array[2244] = 16'h3ece;
mem_array[2247] = 16'h9731;
mem_array[2246] = 16'hbfb2;
mem_array[2249] = 16'h2f36;
mem_array[2248] = 16'hbd94;
mem_array[2251] = 16'h991f;
mem_array[2250] = 16'h3f24;
mem_array[2253] = 16'ha2b6;
mem_array[2252] = 16'h3dcf;
mem_array[2255] = 16'h11dc;
mem_array[2254] = 16'hbe60;
mem_array[2257] = 16'hc763;
mem_array[2256] = 16'h3d7a;
mem_array[2259] = 16'h0c20;
mem_array[2258] = 16'h3edb;
mem_array[2261] = 16'h06a4;
mem_array[2260] = 16'hbd54;
mem_array[2263] = 16'h14bb;
mem_array[2262] = 16'h3e57;
mem_array[2265] = 16'h0c96;
mem_array[2264] = 16'hbe1d;
mem_array[2267] = 16'hfe02;
mem_array[2266] = 16'h3fad;
mem_array[2269] = 16'h9b83;
mem_array[2268] = 16'hbea4;
mem_array[2271] = 16'h330a;
mem_array[2270] = 16'hbde9;
mem_array[2273] = 16'h5e57;
mem_array[2272] = 16'h3e63;
mem_array[2275] = 16'hbbc6;
mem_array[2274] = 16'hbd6f;
mem_array[2277] = 16'h98a0;
mem_array[2276] = 16'hbf3b;
mem_array[2279] = 16'h47a9;
mem_array[2278] = 16'h3db4;
mem_array[2281] = 16'h797a;
mem_array[2280] = 16'hbd02;
mem_array[2283] = 16'he100;
mem_array[2282] = 16'hbd10;
mem_array[2285] = 16'h3210;
mem_array[2284] = 16'h3f20;
mem_array[2287] = 16'h5aca;
mem_array[2286] = 16'h3f66;
mem_array[2289] = 16'h1e3b;
mem_array[2288] = 16'hbe2b;
mem_array[2291] = 16'h6a2b;
mem_array[2290] = 16'h3cc0;
mem_array[2293] = 16'h4982;
mem_array[2292] = 16'hbf42;
mem_array[2295] = 16'h796c;
mem_array[2294] = 16'h3ecf;
mem_array[2297] = 16'h4c1c;
mem_array[2296] = 16'hbf09;
mem_array[2299] = 16'h0ad1;
mem_array[2298] = 16'h3c6c;
mem_array[2301] = 16'h7697;
mem_array[2300] = 16'hbd92;
mem_array[2303] = 16'hc5c4;
mem_array[2302] = 16'h3d39;
mem_array[2305] = 16'habe6;
mem_array[2304] = 16'h3e53;
mem_array[2307] = 16'h7d67;
mem_array[2306] = 16'hbf7d;
mem_array[2309] = 16'hb871;
mem_array[2308] = 16'h3efe;
mem_array[2311] = 16'h4ad3;
mem_array[2310] = 16'h3f23;
mem_array[2313] = 16'hc132;
mem_array[2312] = 16'h3e05;
mem_array[2315] = 16'h1247;
mem_array[2314] = 16'hbe62;
mem_array[2317] = 16'h2162;
mem_array[2316] = 16'h3d9b;
mem_array[2319] = 16'h45aa;
mem_array[2318] = 16'h3efd;
mem_array[2321] = 16'h2696;
mem_array[2320] = 16'hbd93;
mem_array[2323] = 16'h6079;
mem_array[2322] = 16'h3db5;
mem_array[2325] = 16'h9224;
mem_array[2324] = 16'hbd37;
mem_array[2327] = 16'h25fc;
mem_array[2326] = 16'h3fb8;
mem_array[2329] = 16'h7f09;
mem_array[2328] = 16'h3e2f;
mem_array[2331] = 16'h3f6d;
mem_array[2330] = 16'hbd72;
mem_array[2333] = 16'ha588;
mem_array[2332] = 16'h3f1a;
mem_array[2335] = 16'hff53;
mem_array[2334] = 16'h3c9b;
mem_array[2337] = 16'h5591;
mem_array[2336] = 16'hbf23;
mem_array[2339] = 16'hee53;
mem_array[2338] = 16'hbde1;
mem_array[2341] = 16'h4180;
mem_array[2340] = 16'hbc7d;
mem_array[2343] = 16'hb964;
mem_array[2342] = 16'hbd07;
mem_array[2345] = 16'ha59a;
mem_array[2344] = 16'h3ec5;
mem_array[2347] = 16'h9601;
mem_array[2346] = 16'h3e56;
mem_array[2349] = 16'h911e;
mem_array[2348] = 16'hbe8c;
mem_array[2351] = 16'h6887;
mem_array[2350] = 16'hbea2;
mem_array[2353] = 16'hbec8;
mem_array[2352] = 16'hbcd5;
mem_array[2355] = 16'h0fd3;
mem_array[2354] = 16'h3fbb;
mem_array[2357] = 16'h3c61;
mem_array[2356] = 16'hbdff;
mem_array[2359] = 16'hdbf9;
mem_array[2358] = 16'hbf04;
mem_array[2361] = 16'hc0ba;
mem_array[2360] = 16'h3a5d;
mem_array[2363] = 16'hf535;
mem_array[2362] = 16'h3d41;
mem_array[2365] = 16'ha3bd;
mem_array[2364] = 16'h3fc1;
mem_array[2367] = 16'h661c;
mem_array[2366] = 16'hbeda;
mem_array[2369] = 16'hfb64;
mem_array[2368] = 16'h3f24;
mem_array[2371] = 16'hefaf;
mem_array[2370] = 16'hbf98;
mem_array[2373] = 16'hcb95;
mem_array[2372] = 16'h3b0d;
mem_array[2375] = 16'h4be2;
mem_array[2374] = 16'hbf3b;
mem_array[2377] = 16'h7893;
mem_array[2376] = 16'hbe3b;
mem_array[2379] = 16'h4c0d;
mem_array[2378] = 16'hbf82;
mem_array[2381] = 16'h0f89;
mem_array[2380] = 16'hbf50;
mem_array[2383] = 16'h5758;
mem_array[2382] = 16'hbd9f;
mem_array[2385] = 16'h9205;
mem_array[2384] = 16'h3f78;
mem_array[2387] = 16'h238b;
mem_array[2386] = 16'h3f2f;
mem_array[2389] = 16'hb720;
mem_array[2388] = 16'h3e96;
mem_array[2391] = 16'hf473;
mem_array[2390] = 16'hbcdb;
mem_array[2393] = 16'h1a95;
mem_array[2392] = 16'h3f8b;
mem_array[2395] = 16'h3a56;
mem_array[2394] = 16'hbc26;
mem_array[2397] = 16'h2e09;
mem_array[2396] = 16'h3c72;
mem_array[2399] = 16'hb3b6;
mem_array[2398] = 16'hbe9f;
mem_array[2401] = 16'h8b46;
mem_array[2400] = 16'hbcfe;
mem_array[2403] = 16'hf7ed;
mem_array[2402] = 16'h3a2a;
mem_array[2405] = 16'h47a3;
mem_array[2404] = 16'h3e44;
mem_array[2407] = 16'h63e9;
mem_array[2406] = 16'hbd2f;
mem_array[2409] = 16'h2863;
mem_array[2408] = 16'hbd19;
mem_array[2411] = 16'hdf1d;
mem_array[2410] = 16'hbe86;
mem_array[2413] = 16'h31be;
mem_array[2412] = 16'hbe6e;
mem_array[2415] = 16'h7b6e;
mem_array[2414] = 16'h3f64;
mem_array[2417] = 16'hd2eb;
mem_array[2416] = 16'hbe3d;
mem_array[2419] = 16'h3808;
mem_array[2418] = 16'hbea0;
mem_array[2421] = 16'h3164;
mem_array[2420] = 16'h3c69;
mem_array[2423] = 16'h2780;
mem_array[2422] = 16'hbd81;
mem_array[2425] = 16'h5a1f;
mem_array[2424] = 16'h3eca;
mem_array[2427] = 16'h6705;
mem_array[2426] = 16'h3d52;
mem_array[2429] = 16'hbc8a;
mem_array[2428] = 16'h3f12;
mem_array[2431] = 16'h25f4;
mem_array[2430] = 16'hbf12;
mem_array[2433] = 16'h2064;
mem_array[2432] = 16'hbd00;
mem_array[2435] = 16'hd82c;
mem_array[2434] = 16'hbe9f;
mem_array[2437] = 16'h30ce;
mem_array[2436] = 16'hbd24;
mem_array[2439] = 16'h0a98;
mem_array[2438] = 16'hbd9c;
mem_array[2441] = 16'hd3f9;
mem_array[2440] = 16'h3cfe;
mem_array[2443] = 16'hf668;
mem_array[2442] = 16'h3d8f;
mem_array[2445] = 16'h65e6;
mem_array[2444] = 16'h3f50;
mem_array[2447] = 16'h7f44;
mem_array[2446] = 16'h3ef6;
mem_array[2449] = 16'hc9c4;
mem_array[2448] = 16'hbe17;
mem_array[2451] = 16'h13af;
mem_array[2450] = 16'hbd46;
mem_array[2453] = 16'h34af;
mem_array[2452] = 16'h3e01;
mem_array[2455] = 16'hfb5c;
mem_array[2454] = 16'hbd39;
mem_array[2457] = 16'had7c;
mem_array[2456] = 16'hbe3f;
mem_array[2459] = 16'hb4b4;
mem_array[2458] = 16'h3e85;
mem_array[2461] = 16'h9425;
mem_array[2460] = 16'h3d16;
mem_array[2463] = 16'hadc7;
mem_array[2462] = 16'hbce0;
mem_array[2465] = 16'hddc9;
mem_array[2464] = 16'hbe62;
mem_array[2467] = 16'h7cee;
mem_array[2466] = 16'h3e08;
mem_array[2469] = 16'h4f7a;
mem_array[2468] = 16'hbd8e;
mem_array[2471] = 16'h3dd1;
mem_array[2470] = 16'hbf06;
mem_array[2473] = 16'h4b5d;
mem_array[2472] = 16'h3f20;
mem_array[2475] = 16'h0a23;
mem_array[2474] = 16'h3fdc;
mem_array[2477] = 16'hb693;
mem_array[2476] = 16'hbe1e;
mem_array[2479] = 16'h18a1;
mem_array[2478] = 16'h3ea6;
mem_array[2481] = 16'hb77f;
mem_array[2480] = 16'h3d06;
mem_array[2483] = 16'he3f2;
mem_array[2482] = 16'hbcd0;
mem_array[2485] = 16'h5add;
mem_array[2484] = 16'h3f2c;
mem_array[2487] = 16'h2d0a;
mem_array[2486] = 16'hbe14;
mem_array[2489] = 16'h5d3d;
mem_array[2488] = 16'h3e6c;
mem_array[2491] = 16'h4f51;
mem_array[2490] = 16'hbeb7;
mem_array[2493] = 16'hacef;
mem_array[2492] = 16'h3fa1;
mem_array[2495] = 16'h1c54;
mem_array[2494] = 16'hbf7d;
mem_array[2497] = 16'h313e;
mem_array[2496] = 16'hbf23;
mem_array[2499] = 16'h8dde;
mem_array[2498] = 16'h3e48;
mem_array[2501] = 16'h2984;
mem_array[2500] = 16'hbeda;
mem_array[2503] = 16'h8795;
mem_array[2502] = 16'hbe80;
mem_array[2505] = 16'hd598;
mem_array[2504] = 16'h3e80;
mem_array[2507] = 16'hd9ae;
mem_array[2506] = 16'h3ef2;
mem_array[2509] = 16'h8443;
mem_array[2508] = 16'h3cb5;
mem_array[2511] = 16'h0ef8;
mem_array[2510] = 16'hbd14;
mem_array[2513] = 16'h052d;
mem_array[2512] = 16'h3f0a;
mem_array[2515] = 16'ha31c;
mem_array[2514] = 16'hbda3;
mem_array[2517] = 16'hdaca;
mem_array[2516] = 16'h3f5b;
mem_array[2519] = 16'h7e17;
mem_array[2518] = 16'hbda0;
mem_array[2521] = 16'h4373;
mem_array[2520] = 16'hbe3b;
mem_array[2523] = 16'h097c;
mem_array[2522] = 16'hbdf9;
mem_array[2525] = 16'h8b43;
mem_array[2524] = 16'hbe94;
mem_array[2527] = 16'hcef8;
mem_array[2526] = 16'h3e49;
mem_array[2529] = 16'h89a0;
mem_array[2528] = 16'hbd59;
mem_array[2531] = 16'h8329;
mem_array[2530] = 16'hbe06;
mem_array[2533] = 16'h3a13;
mem_array[2532] = 16'hbe7b;
mem_array[2535] = 16'hf5fa;
mem_array[2534] = 16'hbe90;
mem_array[2537] = 16'h7785;
mem_array[2536] = 16'hbcf9;
mem_array[2539] = 16'h318e;
mem_array[2538] = 16'h3e82;
mem_array[2541] = 16'hdbc0;
mem_array[2540] = 16'hbcae;
mem_array[2543] = 16'h1e63;
mem_array[2542] = 16'h3dc7;
mem_array[2545] = 16'h124e;
mem_array[2544] = 16'h3e7f;
mem_array[2547] = 16'hbb93;
mem_array[2546] = 16'hbeee;
mem_array[2549] = 16'h8e87;
mem_array[2548] = 16'hbe26;
mem_array[2551] = 16'hdf20;
mem_array[2550] = 16'hbdf4;
mem_array[2553] = 16'h9f65;
mem_array[2552] = 16'h3f92;
mem_array[2555] = 16'hb5bc;
mem_array[2554] = 16'hbdff;
mem_array[2557] = 16'h317a;
mem_array[2556] = 16'hbe75;
mem_array[2559] = 16'hb306;
mem_array[2558] = 16'hbe63;
mem_array[2561] = 16'heb7a;
mem_array[2560] = 16'hbcc1;
mem_array[2563] = 16'hd6a0;
mem_array[2562] = 16'hbe3b;
mem_array[2565] = 16'heee8;
mem_array[2564] = 16'hbef8;
mem_array[2567] = 16'h28c8;
mem_array[2566] = 16'h3f2c;
mem_array[2569] = 16'h38e1;
mem_array[2568] = 16'hbddb;
mem_array[2571] = 16'h44ad;
mem_array[2570] = 16'h3cc4;
mem_array[2573] = 16'hfed9;
mem_array[2572] = 16'hbe6d;
mem_array[2575] = 16'h5178;
mem_array[2574] = 16'hbd7e;
mem_array[2577] = 16'h1b8f;
mem_array[2576] = 16'hbd5f;
mem_array[2579] = 16'h5e08;
mem_array[2578] = 16'h3f17;
mem_array[2581] = 16'hee4b;
mem_array[2580] = 16'hbec1;
mem_array[2583] = 16'h3000;
mem_array[2582] = 16'hbe8a;
mem_array[2585] = 16'h9df0;
mem_array[2584] = 16'h3e02;
mem_array[2587] = 16'h9e0d;
mem_array[2586] = 16'h3d3d;
mem_array[2589] = 16'hb66c;
mem_array[2588] = 16'hbe5b;
mem_array[2591] = 16'h9bcf;
mem_array[2590] = 16'h3cc7;
mem_array[2593] = 16'hc766;
mem_array[2592] = 16'hbec8;
mem_array[2595] = 16'h5b43;
mem_array[2594] = 16'hbf0b;
mem_array[2597] = 16'h01de;
mem_array[2596] = 16'h3eb8;
mem_array[2599] = 16'hfeb6;
mem_array[2598] = 16'hbe22;
mem_array[2601] = 16'hc3d5;
mem_array[2600] = 16'h3c90;
mem_array[2603] = 16'h01a1;
mem_array[2602] = 16'hbcb5;
mem_array[2605] = 16'h56e0;
mem_array[2604] = 16'h3f3d;
mem_array[2607] = 16'h9e49;
mem_array[2606] = 16'hbe64;
mem_array[2609] = 16'hfbe9;
mem_array[2608] = 16'h3e7d;
mem_array[2611] = 16'h1d97;
mem_array[2610] = 16'hbf03;
mem_array[2613] = 16'hf509;
mem_array[2612] = 16'h3fbd;
mem_array[2615] = 16'had7f;
mem_array[2614] = 16'hbf81;
mem_array[2617] = 16'h36c4;
mem_array[2616] = 16'hbfc8;
mem_array[2619] = 16'h9672;
mem_array[2618] = 16'hbfa4;
mem_array[2621] = 16'h9eee;
mem_array[2620] = 16'hbeb2;
mem_array[2623] = 16'h4118;
mem_array[2622] = 16'h3e26;
mem_array[2625] = 16'h00af;
mem_array[2624] = 16'hbe86;
mem_array[2627] = 16'hee8b;
mem_array[2626] = 16'h3f92;
mem_array[2629] = 16'h1d68;
mem_array[2628] = 16'h3d52;
mem_array[2631] = 16'hf242;
mem_array[2630] = 16'hbea9;
mem_array[2633] = 16'h2d6b;
mem_array[2632] = 16'h3c87;
mem_array[2635] = 16'he0c0;
mem_array[2634] = 16'h3d76;
mem_array[2637] = 16'h89e6;
mem_array[2636] = 16'h3e1b;
mem_array[2639] = 16'h03fe;
mem_array[2638] = 16'h3f0a;
mem_array[2641] = 16'ha451;
mem_array[2640] = 16'hbfc5;
mem_array[2643] = 16'h76fa;
mem_array[2642] = 16'hbdd5;
mem_array[2645] = 16'h01ba;
mem_array[2644] = 16'h3fa3;
mem_array[2647] = 16'he5fd;
mem_array[2646] = 16'h3e4b;
mem_array[2649] = 16'hde95;
mem_array[2648] = 16'h3dfd;
mem_array[2651] = 16'h7b85;
mem_array[2650] = 16'h3d3c;
mem_array[2653] = 16'h945a;
mem_array[2652] = 16'hbf07;
mem_array[2655] = 16'haefe;
mem_array[2654] = 16'hbe41;
mem_array[2657] = 16'h6131;
mem_array[2656] = 16'h3f8d;
mem_array[2659] = 16'hfdd3;
mem_array[2658] = 16'hbf78;
mem_array[2661] = 16'h4ba8;
mem_array[2660] = 16'hbc6b;
mem_array[2663] = 16'hb29a;
mem_array[2662] = 16'h3c4c;
mem_array[2665] = 16'hfe41;
mem_array[2664] = 16'h3ef3;
mem_array[2667] = 16'h6511;
mem_array[2666] = 16'h3f14;
mem_array[2669] = 16'h837d;
mem_array[2668] = 16'h3fb5;
mem_array[2671] = 16'hef7e;
mem_array[2670] = 16'hbf91;
mem_array[2673] = 16'he21d;
mem_array[2672] = 16'h3f7e;
mem_array[2675] = 16'hadef;
mem_array[2674] = 16'hbd91;
mem_array[2677] = 16'h750d;
mem_array[2676] = 16'hbf5d;
mem_array[2679] = 16'h13cf;
mem_array[2678] = 16'hbf99;
mem_array[2681] = 16'h4575;
mem_array[2680] = 16'hbeb4;
mem_array[2683] = 16'hab9f;
mem_array[2682] = 16'h3e9f;
mem_array[2685] = 16'h5f44;
mem_array[2684] = 16'hbf9b;
mem_array[2687] = 16'h28ee;
mem_array[2686] = 16'h3ec7;
mem_array[2689] = 16'h81d1;
mem_array[2688] = 16'h3f26;
mem_array[2691] = 16'hfda5;
mem_array[2690] = 16'h3d82;
mem_array[2693] = 16'h3f85;
mem_array[2692] = 16'h3e28;
mem_array[2695] = 16'h8081;
mem_array[2694] = 16'h3d4a;
mem_array[2697] = 16'h423e;
mem_array[2696] = 16'h3f86;
mem_array[2699] = 16'hf2f8;
mem_array[2698] = 16'hbe5a;
mem_array[2701] = 16'h2fb9;
mem_array[2700] = 16'hbe97;
mem_array[2703] = 16'h4296;
mem_array[2702] = 16'hbcf4;
mem_array[2705] = 16'h2f92;
mem_array[2704] = 16'h3f64;
mem_array[2707] = 16'he8c3;
mem_array[2706] = 16'h3e52;
mem_array[2709] = 16'h530d;
mem_array[2708] = 16'h3e80;
mem_array[2711] = 16'h82e0;
mem_array[2710] = 16'h3e22;
mem_array[2713] = 16'h8525;
mem_array[2712] = 16'hbe1e;
mem_array[2715] = 16'h3165;
mem_array[2714] = 16'h3e89;
mem_array[2717] = 16'h6f30;
mem_array[2716] = 16'h3de9;
mem_array[2719] = 16'h1253;
mem_array[2718] = 16'hbe11;
mem_array[2721] = 16'h4e07;
mem_array[2720] = 16'hbdc2;
mem_array[2723] = 16'hdf5a;
mem_array[2722] = 16'hbda1;
mem_array[2725] = 16'h37e6;
mem_array[2724] = 16'h3f7a;
mem_array[2727] = 16'h73d2;
mem_array[2726] = 16'hbc58;
mem_array[2729] = 16'h1e2a;
mem_array[2728] = 16'h3ebf;
mem_array[2731] = 16'h4356;
mem_array[2730] = 16'hbf54;
mem_array[2733] = 16'h9f28;
mem_array[2732] = 16'h3f62;
mem_array[2735] = 16'hb186;
mem_array[2734] = 16'hbdc8;
mem_array[2737] = 16'h9ac7;
mem_array[2736] = 16'hbd98;
mem_array[2739] = 16'h5b77;
mem_array[2738] = 16'hbf8a;
mem_array[2741] = 16'h08ce;
mem_array[2740] = 16'hbe5b;
mem_array[2743] = 16'h2a89;
mem_array[2742] = 16'h3e00;
mem_array[2745] = 16'h65ea;
mem_array[2744] = 16'h3ea6;
mem_array[2747] = 16'ha7e8;
mem_array[2746] = 16'h3ecf;
mem_array[2749] = 16'hc362;
mem_array[2748] = 16'hbe26;
mem_array[2751] = 16'hee9d;
mem_array[2750] = 16'hbbf2;
mem_array[2753] = 16'hc58d;
mem_array[2752] = 16'h3e0f;
mem_array[2755] = 16'hcd42;
mem_array[2754] = 16'h3b8a;
mem_array[2757] = 16'hd6e7;
mem_array[2756] = 16'hbe67;
mem_array[2759] = 16'h807a;
mem_array[2758] = 16'h3e03;
mem_array[2761] = 16'h1c95;
mem_array[2760] = 16'h3d83;
mem_array[2763] = 16'hacd0;
mem_array[2762] = 16'h3c04;
mem_array[2765] = 16'h9753;
mem_array[2764] = 16'h3e37;
mem_array[2767] = 16'hf7ff;
mem_array[2766] = 16'hbea3;
mem_array[2769] = 16'h32ae;
mem_array[2768] = 16'hbd8d;
mem_array[2771] = 16'h26e3;
mem_array[2770] = 16'h3d23;
mem_array[2773] = 16'hfcbe;
mem_array[2772] = 16'hbd90;
mem_array[2775] = 16'h7ae9;
mem_array[2774] = 16'h3e8e;
mem_array[2777] = 16'h0c12;
mem_array[2776] = 16'hbe55;
mem_array[2779] = 16'hb2ce;
mem_array[2778] = 16'hbf36;
mem_array[2781] = 16'h1962;
mem_array[2780] = 16'hbd09;
mem_array[2783] = 16'h8c51;
mem_array[2782] = 16'hb987;
mem_array[2785] = 16'h2441;
mem_array[2784] = 16'h3f90;
mem_array[2787] = 16'hd20c;
mem_array[2786] = 16'hbe14;
mem_array[2789] = 16'h2205;
mem_array[2788] = 16'hbe32;
mem_array[2791] = 16'hbe2c;
mem_array[2790] = 16'hbfda;
mem_array[2793] = 16'hbfb4;
mem_array[2792] = 16'h3ef9;
mem_array[2795] = 16'h9dfb;
mem_array[2794] = 16'h3dcc;
mem_array[2797] = 16'h8d2d;
mem_array[2796] = 16'h3ddf;
mem_array[2799] = 16'h2c72;
mem_array[2798] = 16'hbf0e;
mem_array[2801] = 16'h159a;
mem_array[2800] = 16'hbe7e;
mem_array[2803] = 16'hfd91;
mem_array[2802] = 16'hbeaf;
mem_array[2805] = 16'hc702;
mem_array[2804] = 16'h3f94;
mem_array[2807] = 16'he808;
mem_array[2806] = 16'h3f09;
mem_array[2809] = 16'h932b;
mem_array[2808] = 16'hbdc1;
mem_array[2811] = 16'h0f9a;
mem_array[2810] = 16'hbd7d;
mem_array[2813] = 16'hc6c7;
mem_array[2812] = 16'hbeef;
mem_array[2815] = 16'hc0b1;
mem_array[2814] = 16'h3f52;
mem_array[2817] = 16'hf5ae;
mem_array[2816] = 16'hbe63;
mem_array[2819] = 16'h0475;
mem_array[2818] = 16'hbcee;
mem_array[2821] = 16'h0e69;
mem_array[2820] = 16'h3d5c;
mem_array[2823] = 16'h418d;
mem_array[2822] = 16'hbc54;
mem_array[2825] = 16'h47fc;
mem_array[2824] = 16'h3cbb;
mem_array[2827] = 16'h438d;
mem_array[2826] = 16'h3d9c;
mem_array[2829] = 16'hcc3e;
mem_array[2828] = 16'h3d2b;
mem_array[2831] = 16'h9704;
mem_array[2830] = 16'h3e86;
mem_array[2833] = 16'h4e2a;
mem_array[2832] = 16'hbeef;
mem_array[2835] = 16'h202a;
mem_array[2834] = 16'hbe42;
mem_array[2837] = 16'h48f1;
mem_array[2836] = 16'h3f1e;
mem_array[2839] = 16'h6092;
mem_array[2838] = 16'h3d02;
mem_array[2841] = 16'h621c;
mem_array[2840] = 16'h3dcf;
mem_array[2843] = 16'h3d72;
mem_array[2842] = 16'hbd22;
mem_array[2845] = 16'h96a9;
mem_array[2844] = 16'h3f56;
mem_array[2847] = 16'hc83b;
mem_array[2846] = 16'h3d42;
mem_array[2849] = 16'hf061;
mem_array[2848] = 16'h3d9c;
mem_array[2851] = 16'h3c17;
mem_array[2850] = 16'hbdde;
mem_array[2853] = 16'h72ce;
mem_array[2852] = 16'hbd45;
mem_array[2855] = 16'h5f70;
mem_array[2854] = 16'h3cef;
mem_array[2857] = 16'h5a12;
mem_array[2856] = 16'hbf0f;
mem_array[2859] = 16'hd315;
mem_array[2858] = 16'h3ee9;
mem_array[2861] = 16'h1dac;
mem_array[2860] = 16'hbdce;
mem_array[2863] = 16'h2246;
mem_array[2862] = 16'hbe0c;
mem_array[2865] = 16'h974c;
mem_array[2864] = 16'hbe91;
mem_array[2867] = 16'h9fd5;
mem_array[2866] = 16'h3a8a;
mem_array[2869] = 16'hcc95;
mem_array[2868] = 16'h3d0a;
mem_array[2871] = 16'h766e;
mem_array[2870] = 16'h3d7b;
mem_array[2873] = 16'h2e36;
mem_array[2872] = 16'hbdbc;
mem_array[2875] = 16'h8e49;
mem_array[2874] = 16'h3d2d;
mem_array[2877] = 16'h5c35;
mem_array[2876] = 16'hbda7;
mem_array[2879] = 16'h7526;
mem_array[2878] = 16'h3de6;
mem_array[2881] = 16'h1e14;
mem_array[2880] = 16'hbc9e;
mem_array[2883] = 16'hc621;
mem_array[2882] = 16'hbc3a;
mem_array[2885] = 16'h5d1c;
mem_array[2884] = 16'h3c23;
mem_array[2887] = 16'h5a7e;
mem_array[2886] = 16'h3c68;
mem_array[2889] = 16'h57c0;
mem_array[2888] = 16'hbc88;
mem_array[2891] = 16'h6c7d;
mem_array[2890] = 16'h3ea0;
mem_array[2893] = 16'h396e;
mem_array[2892] = 16'hbd9a;
mem_array[2895] = 16'h1e70;
mem_array[2894] = 16'hbdf2;
mem_array[2897] = 16'h03b6;
mem_array[2896] = 16'h3f0b;
mem_array[2899] = 16'h0b3f;
mem_array[2898] = 16'hbd13;
mem_array[2901] = 16'hb382;
mem_array[2900] = 16'h3e11;
mem_array[2903] = 16'h1b70;
mem_array[2902] = 16'hbd44;
mem_array[2905] = 16'h4eef;
mem_array[2904] = 16'h3f53;
mem_array[2907] = 16'h380c;
mem_array[2906] = 16'h3c4c;
mem_array[2909] = 16'h004a;
mem_array[2908] = 16'hbd99;
mem_array[2911] = 16'h95ad;
mem_array[2910] = 16'hbe8e;
mem_array[2913] = 16'h96d3;
mem_array[2912] = 16'hbce2;
mem_array[2915] = 16'hd826;
mem_array[2914] = 16'hbde7;
mem_array[2917] = 16'h74fb;
mem_array[2916] = 16'hbeca;
mem_array[2919] = 16'hdc13;
mem_array[2918] = 16'hbed3;
mem_array[2921] = 16'hd6f1;
mem_array[2920] = 16'hbe4e;
mem_array[2923] = 16'h3702;
mem_array[2922] = 16'h3d3c;
mem_array[2925] = 16'h9b2e;
mem_array[2924] = 16'h3ecd;
mem_array[2927] = 16'hfaeb;
mem_array[2926] = 16'h3e87;
mem_array[2929] = 16'hd295;
mem_array[2928] = 16'h3a90;
mem_array[2931] = 16'hd00f;
mem_array[2930] = 16'hbd2c;
mem_array[2933] = 16'hd9a1;
mem_array[2932] = 16'h3d51;
mem_array[2935] = 16'h4749;
mem_array[2934] = 16'hbd6e;
mem_array[2937] = 16'h398a;
mem_array[2936] = 16'hbd62;
mem_array[2939] = 16'h8f7f;
mem_array[2938] = 16'hbb18;
mem_array[2941] = 16'h3022;
mem_array[2940] = 16'h3da4;
mem_array[2943] = 16'h1107;
mem_array[2942] = 16'h3db1;
mem_array[2945] = 16'hc542;
mem_array[2944] = 16'hbc22;
mem_array[2947] = 16'he9de;
mem_array[2946] = 16'hbc14;
mem_array[2949] = 16'h38f9;
mem_array[2948] = 16'hbce7;
mem_array[2951] = 16'h0435;
mem_array[2950] = 16'h3ee5;
mem_array[2953] = 16'h336b;
mem_array[2952] = 16'hbeca;
mem_array[2955] = 16'h48b2;
mem_array[2954] = 16'hbe4b;
mem_array[2957] = 16'hd138;
mem_array[2956] = 16'hbd97;
mem_array[2959] = 16'h2e85;
mem_array[2958] = 16'h3c0f;
mem_array[2961] = 16'h3ce8;
mem_array[2960] = 16'h3cef;
mem_array[2963] = 16'hc2f7;
mem_array[2962] = 16'hbc13;
mem_array[2965] = 16'h6d55;
mem_array[2964] = 16'h3f27;
mem_array[2967] = 16'h3f7b;
mem_array[2966] = 16'hbe28;
mem_array[2969] = 16'h544b;
mem_array[2968] = 16'hbe40;
mem_array[2971] = 16'h8ac9;
mem_array[2970] = 16'hbc8c;
mem_array[2973] = 16'h987d;
mem_array[2972] = 16'h3d6f;
mem_array[2975] = 16'hb86c;
mem_array[2974] = 16'hbd9e;
mem_array[2977] = 16'hd094;
mem_array[2976] = 16'hbe41;
mem_array[2979] = 16'h8c36;
mem_array[2978] = 16'h3e13;
mem_array[2981] = 16'h0f6b;
mem_array[2980] = 16'hbd5b;
mem_array[2983] = 16'h75b4;
mem_array[2982] = 16'h3e05;
mem_array[2985] = 16'hd756;
mem_array[2984] = 16'h3e40;
mem_array[2987] = 16'ha13f;
mem_array[2986] = 16'h3d1b;
mem_array[2989] = 16'hcc60;
mem_array[2988] = 16'h3dec;
mem_array[2991] = 16'h48a5;
mem_array[2990] = 16'hba27;
mem_array[2993] = 16'h1661;
mem_array[2992] = 16'hbe40;
mem_array[2995] = 16'h8dc0;
mem_array[2994] = 16'h3cb3;
mem_array[2997] = 16'hb015;
mem_array[2996] = 16'hbc5a;
mem_array[2999] = 16'he069;
mem_array[2998] = 16'hbce1;
mem_array[3001] = 16'hcfde;
mem_array[3000] = 16'h3d84;
mem_array[3003] = 16'h4051;
mem_array[3002] = 16'h3d19;
mem_array[3005] = 16'h70f5;
mem_array[3004] = 16'h3dc6;
mem_array[3007] = 16'he4f5;
mem_array[3006] = 16'hbbb4;
mem_array[3009] = 16'hb35e;
mem_array[3008] = 16'hbe0a;
mem_array[3011] = 16'hf361;
mem_array[3010] = 16'h3ec9;
mem_array[3013] = 16'h46c4;
mem_array[3012] = 16'hbe8b;
mem_array[3015] = 16'h8f00;
mem_array[3014] = 16'hbec7;
mem_array[3017] = 16'hb9f8;
mem_array[3016] = 16'hbe79;
mem_array[3019] = 16'h5956;
mem_array[3018] = 16'h3e01;
mem_array[3021] = 16'heef6;
mem_array[3020] = 16'h3d99;
mem_array[3023] = 16'h0d26;
mem_array[3022] = 16'hbddb;
mem_array[3025] = 16'h7290;
mem_array[3024] = 16'h3f61;
mem_array[3027] = 16'hba36;
mem_array[3026] = 16'h3d0a;
mem_array[3029] = 16'h6c60;
mem_array[3028] = 16'hbe42;
mem_array[3031] = 16'ha358;
mem_array[3030] = 16'h3d41;
mem_array[3033] = 16'hb836;
mem_array[3032] = 16'h3d88;
mem_array[3035] = 16'hb80b;
mem_array[3034] = 16'hbd06;
mem_array[3037] = 16'h9ce7;
mem_array[3036] = 16'hbe8f;
mem_array[3039] = 16'h9ce1;
mem_array[3038] = 16'h3e72;
mem_array[3041] = 16'h72f1;
mem_array[3040] = 16'hbdbf;
mem_array[3043] = 16'hcac3;
mem_array[3042] = 16'h3d04;
mem_array[3045] = 16'h1eb7;
mem_array[3044] = 16'h3ded;
mem_array[3047] = 16'h74bc;
mem_array[3046] = 16'h3e2e;
mem_array[3049] = 16'hd846;
mem_array[3048] = 16'h3e8a;
mem_array[3051] = 16'h1597;
mem_array[3050] = 16'hbd0d;
mem_array[3053] = 16'h97ed;
mem_array[3052] = 16'hbe46;
mem_array[3055] = 16'haed2;
mem_array[3054] = 16'hbda2;
mem_array[3057] = 16'hbebf;
mem_array[3056] = 16'hbd47;
mem_array[3059] = 16'ha611;
mem_array[3058] = 16'hbe3b;
mem_array[3061] = 16'hc76d;
mem_array[3060] = 16'hbd5f;
mem_array[3063] = 16'hb2c4;
mem_array[3062] = 16'h3d6f;
mem_array[3065] = 16'hfc5f;
mem_array[3064] = 16'hbb90;
mem_array[3067] = 16'h87cb;
mem_array[3066] = 16'h3d9b;
mem_array[3069] = 16'hf19e;
mem_array[3068] = 16'h3cc8;
mem_array[3071] = 16'h8372;
mem_array[3070] = 16'hbd93;
mem_array[3073] = 16'hdd60;
mem_array[3072] = 16'hbd15;
mem_array[3075] = 16'hded6;
mem_array[3074] = 16'h3ce0;
mem_array[3077] = 16'h2fa2;
mem_array[3076] = 16'hbd86;
mem_array[3079] = 16'hd264;
mem_array[3078] = 16'hbc89;
mem_array[3081] = 16'h6f48;
mem_array[3080] = 16'hbde3;
mem_array[3083] = 16'h6e7d;
mem_array[3082] = 16'h3d10;
mem_array[3085] = 16'hd0f0;
mem_array[3084] = 16'h3e07;
mem_array[3087] = 16'h663b;
mem_array[3086] = 16'hbd4e;
mem_array[3089] = 16'h4338;
mem_array[3088] = 16'h3d18;
mem_array[3091] = 16'h01dc;
mem_array[3090] = 16'hbd9b;
mem_array[3093] = 16'he375;
mem_array[3092] = 16'h3cc1;
mem_array[3095] = 16'hd5fa;
mem_array[3094] = 16'hbded;
mem_array[3097] = 16'h6f74;
mem_array[3096] = 16'hbdc8;
mem_array[3099] = 16'h3ea9;
mem_array[3098] = 16'hbd0f;
mem_array[3101] = 16'hb54a;
mem_array[3100] = 16'hbe17;
mem_array[3103] = 16'h63e5;
mem_array[3102] = 16'h3dd1;
mem_array[3105] = 16'h5700;
mem_array[3104] = 16'hbcdf;
mem_array[3107] = 16'h00bd;
mem_array[3106] = 16'h3d0f;
mem_array[3109] = 16'h2cc5;
mem_array[3108] = 16'h3c80;
mem_array[3111] = 16'h8496;
mem_array[3110] = 16'h3c90;
mem_array[3113] = 16'h8eee;
mem_array[3112] = 16'h3d3d;
mem_array[3115] = 16'h86b7;
mem_array[3114] = 16'hbbc4;
mem_array[3117] = 16'hf6b3;
mem_array[3116] = 16'hbcc7;
mem_array[3119] = 16'h39bf;
mem_array[3118] = 16'hbd34;
mem_array[3121] = 16'h4d6e;
mem_array[3120] = 16'hbd46;
mem_array[3123] = 16'h02d5;
mem_array[3122] = 16'h3ba2;
mem_array[3125] = 16'h1771;
mem_array[3124] = 16'h3dc1;
mem_array[3127] = 16'he00a;
mem_array[3126] = 16'h3d81;
mem_array[3129] = 16'h072a;
mem_array[3128] = 16'hbc47;
mem_array[3131] = 16'hd909;
mem_array[3130] = 16'h3c95;
mem_array[3133] = 16'h9c07;
mem_array[3132] = 16'h3c60;
mem_array[3135] = 16'h14f6;
mem_array[3134] = 16'h3d1d;
mem_array[3137] = 16'h51a2;
mem_array[3136] = 16'hbc9d;
mem_array[3139] = 16'h5157;
mem_array[3138] = 16'h3d80;
mem_array[3141] = 16'h6d09;
mem_array[3140] = 16'h3dc4;
mem_array[3143] = 16'h8719;
mem_array[3142] = 16'hbd3c;
mem_array[3145] = 16'h49db;
mem_array[3144] = 16'hbd7c;
mem_array[3147] = 16'hab23;
mem_array[3146] = 16'hbc2c;
mem_array[3149] = 16'h6cf7;
mem_array[3148] = 16'hbdb6;
mem_array[3151] = 16'hf892;
mem_array[3150] = 16'hbd44;
mem_array[3153] = 16'hb4e3;
mem_array[3152] = 16'hbcc4;
mem_array[3155] = 16'h3d3b;
mem_array[3154] = 16'h3d26;
mem_array[3157] = 16'h39a7;
mem_array[3156] = 16'h3c1c;
mem_array[3159] = 16'hbaad;
mem_array[3158] = 16'h3c94;
mem_array[3161] = 16'hc499;
mem_array[3160] = 16'h3c9f;
mem_array[3163] = 16'ha731;
mem_array[3162] = 16'hbcc0;
mem_array[3165] = 16'h1ae6;
mem_array[3164] = 16'h3d6c;
mem_array[3167] = 16'h2d32;
mem_array[3166] = 16'hbd8b;
mem_array[3169] = 16'h3c82;
mem_array[3168] = 16'hbb05;
mem_array[3171] = 16'hf5d3;
mem_array[3170] = 16'h3c7b;
mem_array[3173] = 16'hbd38;
mem_array[3172] = 16'h3d7a;
mem_array[3175] = 16'ha69a;
mem_array[3174] = 16'hbdb8;
mem_array[3177] = 16'h9660;
mem_array[3176] = 16'hbc95;
mem_array[3179] = 16'h68be;
mem_array[3178] = 16'hbd88;
mem_array[3181] = 16'hc4a0;
mem_array[3180] = 16'h3cb3;
mem_array[3183] = 16'h4f19;
mem_array[3182] = 16'h3cdc;
mem_array[3185] = 16'hb110;
mem_array[3184] = 16'h3d78;
mem_array[3187] = 16'hc1e9;
mem_array[3186] = 16'h3cd6;
mem_array[3189] = 16'h4b5d;
mem_array[3188] = 16'hbd2f;
mem_array[3191] = 16'he9b9;
mem_array[3190] = 16'hbd06;
mem_array[3193] = 16'hee71;
mem_array[3192] = 16'hbc74;
mem_array[3195] = 16'h5e81;
mem_array[3194] = 16'hbd8a;
mem_array[3197] = 16'hf487;
mem_array[3196] = 16'h3cff;
mem_array[3199] = 16'hf591;
mem_array[3198] = 16'h3d56;
mem_array[3201] = 16'h5ac1;
mem_array[3200] = 16'h3dd9;
mem_array[3203] = 16'h2606;
mem_array[3202] = 16'h3cd7;
mem_array[3205] = 16'h9554;
mem_array[3204] = 16'h3d24;
mem_array[3207] = 16'hd851;
mem_array[3206] = 16'h3c57;
mem_array[3209] = 16'hf9be;
mem_array[3208] = 16'hbd02;
mem_array[3211] = 16'hf4e1;
mem_array[3210] = 16'h3d16;
mem_array[3213] = 16'haff5;
mem_array[3212] = 16'hbde9;
mem_array[3215] = 16'h33fb;
mem_array[3214] = 16'h3d97;
mem_array[3217] = 16'h7e70;
mem_array[3216] = 16'h3d96;
mem_array[3219] = 16'h2a51;
mem_array[3218] = 16'hbd5a;
mem_array[3221] = 16'hbebd;
mem_array[3220] = 16'h3c90;
mem_array[3223] = 16'h0bf0;
mem_array[3222] = 16'hbcb5;
mem_array[3225] = 16'h9d40;
mem_array[3224] = 16'hbba8;
mem_array[3227] = 16'heb09;
mem_array[3226] = 16'hbcc2;
mem_array[3229] = 16'h693b;
mem_array[3228] = 16'hbdbc;
mem_array[3231] = 16'h9c44;
mem_array[3230] = 16'hbc1e;
mem_array[3233] = 16'h4405;
mem_array[3232] = 16'h3cbb;
mem_array[3235] = 16'hc262;
mem_array[3234] = 16'h3da2;
mem_array[3237] = 16'hb4bb;
mem_array[3236] = 16'hbd17;
mem_array[3239] = 16'h22e5;
mem_array[3238] = 16'hbd34;
mem_array[3241] = 16'h1894;
mem_array[3240] = 16'h3d15;
mem_array[3243] = 16'hf7de;
mem_array[3242] = 16'h3d89;
mem_array[3245] = 16'h8861;
mem_array[3244] = 16'h3dc6;
mem_array[3247] = 16'h221f;
mem_array[3246] = 16'h3c74;
mem_array[3249] = 16'hf82c;
mem_array[3248] = 16'h3c5d;
mem_array[3251] = 16'he35b;
mem_array[3250] = 16'h3d2d;
mem_array[3253] = 16'h39b2;
mem_array[3252] = 16'hbc51;
mem_array[3255] = 16'h342c;
mem_array[3254] = 16'h3d15;
mem_array[3257] = 16'hf14c;
mem_array[3256] = 16'hbdb8;
mem_array[3259] = 16'ha105;
mem_array[3258] = 16'hbd73;
mem_array[3261] = 16'h238f;
mem_array[3260] = 16'hbd83;
mem_array[3263] = 16'hc580;
mem_array[3262] = 16'hbcb5;
mem_array[3265] = 16'ha97c;
mem_array[3264] = 16'hbd97;
mem_array[3267] = 16'hd2dc;
mem_array[3266] = 16'hbce9;
mem_array[3269] = 16'h54cc;
mem_array[3268] = 16'hbd88;
mem_array[3271] = 16'h9450;
mem_array[3270] = 16'hbcef;
mem_array[3273] = 16'hf6bd;
mem_array[3272] = 16'hbc41;
mem_array[3275] = 16'h8e47;
mem_array[3274] = 16'hbd04;
mem_array[3277] = 16'h561c;
mem_array[3276] = 16'hbdc6;
mem_array[3279] = 16'hfafe;
mem_array[3278] = 16'h3da2;
mem_array[3281] = 16'h592b;
mem_array[3280] = 16'hbbe4;
mem_array[3283] = 16'hddf8;
mem_array[3282] = 16'h3bb6;
mem_array[3285] = 16'h7857;
mem_array[3284] = 16'h3db1;
mem_array[3287] = 16'h7dc1;
mem_array[3286] = 16'hbd4f;
mem_array[3289] = 16'h76ff;
mem_array[3288] = 16'h3db0;
mem_array[3291] = 16'h80ba;
mem_array[3290] = 16'h3ca2;
mem_array[3293] = 16'h0beb;
mem_array[3292] = 16'h3ae9;
mem_array[3295] = 16'h1f37;
mem_array[3294] = 16'hbd06;
mem_array[3297] = 16'h46bc;
mem_array[3296] = 16'h3da3;
mem_array[3299] = 16'hc136;
mem_array[3298] = 16'h3d08;
mem_array[3301] = 16'hcf1e;
mem_array[3300] = 16'hbb59;
mem_array[3303] = 16'h647f;
mem_array[3302] = 16'hbd07;
mem_array[3305] = 16'hf0f0;
mem_array[3304] = 16'h3d2c;
mem_array[3307] = 16'h8e3d;
mem_array[3306] = 16'hba3c;
mem_array[3309] = 16'h4005;
mem_array[3308] = 16'h3cc7;
mem_array[3311] = 16'ha083;
mem_array[3310] = 16'h3d24;
mem_array[3313] = 16'hb26c;
mem_array[3312] = 16'hba1c;
mem_array[3315] = 16'h60c8;
mem_array[3314] = 16'h3d39;
mem_array[3317] = 16'hb225;
mem_array[3316] = 16'hbd14;
mem_array[3319] = 16'h584e;
mem_array[3318] = 16'hbd47;
mem_array[3321] = 16'h2ef6;
mem_array[3320] = 16'h3da7;
mem_array[3323] = 16'h6ac9;
mem_array[3322] = 16'hbc3d;
mem_array[3325] = 16'h9520;
mem_array[3324] = 16'hbce7;
mem_array[3327] = 16'h307b;
mem_array[3326] = 16'hbce4;
mem_array[3329] = 16'h13bd;
mem_array[3328] = 16'h3d7f;
mem_array[3331] = 16'h6fdb;
mem_array[3330] = 16'h3cee;
mem_array[3333] = 16'h4285;
mem_array[3332] = 16'hbbe3;
mem_array[3335] = 16'h7999;
mem_array[3334] = 16'hbd0e;
mem_array[3337] = 16'had3d;
mem_array[3336] = 16'hbb96;
mem_array[3339] = 16'h1275;
mem_array[3338] = 16'h3d9c;
mem_array[3341] = 16'hfd7c;
mem_array[3340] = 16'hbbd4;
mem_array[3343] = 16'h2e59;
mem_array[3342] = 16'hbca1;
mem_array[3345] = 16'h28ac;
mem_array[3344] = 16'h3d52;
mem_array[3347] = 16'h62ae;
mem_array[3346] = 16'hbce8;
mem_array[3349] = 16'h4c89;
mem_array[3348] = 16'hbca5;
mem_array[3351] = 16'h27af;
mem_array[3350] = 16'hbb9c;
mem_array[3353] = 16'h63ca;
mem_array[3352] = 16'hbcd5;
mem_array[3355] = 16'h7712;
mem_array[3354] = 16'h3da8;
mem_array[3357] = 16'h9588;
mem_array[3356] = 16'hbd73;
mem_array[3359] = 16'h3387;
mem_array[3358] = 16'hbba0;
mem_array[3361] = 16'h6843;
mem_array[3360] = 16'h3c86;
mem_array[3363] = 16'h22cd;
mem_array[3362] = 16'h3dbc;
mem_array[3365] = 16'h8a29;
mem_array[3364] = 16'hbd25;
mem_array[3367] = 16'hf940;
mem_array[3366] = 16'hbd43;
mem_array[3369] = 16'h9ea2;
mem_array[3368] = 16'hbd80;
mem_array[3371] = 16'hc2c1;
mem_array[3370] = 16'h3d70;
mem_array[3373] = 16'haac6;
mem_array[3372] = 16'h3ac7;
mem_array[3375] = 16'h1ffe;
mem_array[3374] = 16'hbd18;
mem_array[3377] = 16'h1327;
mem_array[3376] = 16'h3d2d;
mem_array[3379] = 16'h7c78;
mem_array[3378] = 16'h3d9a;
mem_array[3381] = 16'h04cf;
mem_array[3380] = 16'hbc82;
mem_array[3383] = 16'hccf4;
mem_array[3382] = 16'hbd5d;
mem_array[3385] = 16'h3043;
mem_array[3384] = 16'h3d7a;
mem_array[3387] = 16'hc1c7;
mem_array[3386] = 16'hbcdb;
mem_array[3389] = 16'h7959;
mem_array[3388] = 16'hbc5b;
mem_array[3391] = 16'h1039;
mem_array[3390] = 16'hbd19;
mem_array[3393] = 16'hf464;
mem_array[3392] = 16'hbd5c;
mem_array[3395] = 16'h7a60;
mem_array[3394] = 16'h3c4e;
mem_array[3397] = 16'hbc14;
mem_array[3396] = 16'h3b3d;
mem_array[3399] = 16'hd58b;
mem_array[3398] = 16'hbc10;
mem_array[3401] = 16'hb862;
mem_array[3400] = 16'hbdb8;
mem_array[3403] = 16'hf8e4;
mem_array[3402] = 16'hbde5;
mem_array[3405] = 16'h6c6e;
mem_array[3404] = 16'h3cf7;
mem_array[3407] = 16'h7abc;
mem_array[3406] = 16'h3d21;
mem_array[3409] = 16'h4274;
mem_array[3408] = 16'hbde4;
mem_array[3411] = 16'h8561;
mem_array[3410] = 16'h3d1b;
mem_array[3413] = 16'h3524;
mem_array[3412] = 16'h3d23;
mem_array[3415] = 16'hf9f4;
mem_array[3414] = 16'h3d90;
mem_array[3417] = 16'h3db9;
mem_array[3416] = 16'hbc61;
mem_array[3419] = 16'h729e;
mem_array[3418] = 16'hbd85;
mem_array[3421] = 16'hcc03;
mem_array[3420] = 16'hbc7c;
mem_array[3423] = 16'h2367;
mem_array[3422] = 16'hbd19;
mem_array[3425] = 16'h7dfd;
mem_array[3424] = 16'h3d04;
mem_array[3427] = 16'h48c8;
mem_array[3426] = 16'h3c49;
mem_array[3429] = 16'h6175;
mem_array[3428] = 16'h3d7c;
mem_array[3431] = 16'h4ce0;
mem_array[3430] = 16'hbd08;
mem_array[3433] = 16'h787a;
mem_array[3432] = 16'h3c4c;
mem_array[3435] = 16'h4aa0;
mem_array[3434] = 16'h3c8e;
mem_array[3437] = 16'h131c;
mem_array[3436] = 16'h3d6a;
mem_array[3439] = 16'hc44f;
mem_array[3438] = 16'h3dac;
mem_array[3441] = 16'haec2;
mem_array[3440] = 16'hbc6d;
mem_array[3443] = 16'h0def;
mem_array[3442] = 16'hbd22;
mem_array[3445] = 16'h8f0e;
mem_array[3444] = 16'hbcf0;
mem_array[3447] = 16'hd35b;
mem_array[3446] = 16'h3cff;
mem_array[3449] = 16'haa84;
mem_array[3448] = 16'h3d30;
mem_array[3451] = 16'hba51;
mem_array[3450] = 16'h3d3d;
mem_array[3453] = 16'h7790;
mem_array[3452] = 16'h3bd0;
mem_array[3455] = 16'he665;
mem_array[3454] = 16'hbd1f;
mem_array[3457] = 16'h5900;
mem_array[3456] = 16'hbdb3;
mem_array[3459] = 16'h0c0a;
mem_array[3458] = 16'hbd8f;
mem_array[3461] = 16'h5ae8;
mem_array[3460] = 16'h3db7;
mem_array[3463] = 16'h64c0;
mem_array[3462] = 16'hbd30;
mem_array[3465] = 16'hd22d;
mem_array[3464] = 16'hbdaf;
mem_array[3467] = 16'h2f33;
mem_array[3466] = 16'hbd51;
mem_array[3469] = 16'h2f2d;
mem_array[3468] = 16'hb992;
mem_array[3471] = 16'h6483;
mem_array[3470] = 16'h3b31;
mem_array[3473] = 16'h5a0d;
mem_array[3472] = 16'hbd7b;
mem_array[3475] = 16'h0963;
mem_array[3474] = 16'h3cdc;
mem_array[3477] = 16'hb5ab;
mem_array[3476] = 16'hbd79;
mem_array[3479] = 16'hed86;
mem_array[3478] = 16'hbcea;
mem_array[3481] = 16'h87d5;
mem_array[3480] = 16'hbd8d;
mem_array[3483] = 16'h434c;
mem_array[3482] = 16'hbcbf;
mem_array[3485] = 16'h57d1;
mem_array[3484] = 16'h3c8f;
mem_array[3487] = 16'hf598;
mem_array[3486] = 16'h3d0a;
mem_array[3489] = 16'h3b52;
mem_array[3488] = 16'hbbe0;
mem_array[3491] = 16'h33d0;
mem_array[3490] = 16'hbccd;
mem_array[3493] = 16'h6312;
mem_array[3492] = 16'h3c9e;
mem_array[3495] = 16'hcbe3;
mem_array[3494] = 16'h3d17;
mem_array[3497] = 16'h6308;
mem_array[3496] = 16'hbcfe;
mem_array[3499] = 16'hb785;
mem_array[3498] = 16'h3d98;
mem_array[3501] = 16'h9511;
mem_array[3500] = 16'h3dba;
mem_array[3503] = 16'h11fb;
mem_array[3502] = 16'h3c44;
mem_array[3505] = 16'h66f2;
mem_array[3504] = 16'h3ce6;
mem_array[3507] = 16'haba2;
mem_array[3506] = 16'h3ce4;
mem_array[3509] = 16'h4d88;
mem_array[3508] = 16'h3d96;
mem_array[3511] = 16'hffe2;
mem_array[3510] = 16'h3af9;
mem_array[3513] = 16'hbf8f;
mem_array[3512] = 16'h3ce3;
mem_array[3515] = 16'h4cac;
mem_array[3514] = 16'hbb85;
mem_array[3517] = 16'h5661;
mem_array[3516] = 16'hbd90;
mem_array[3519] = 16'hf96f;
mem_array[3518] = 16'h3d91;
mem_array[3521] = 16'hb4ab;
mem_array[3520] = 16'hbdde;
mem_array[3523] = 16'h455e;
mem_array[3522] = 16'h3d5b;
mem_array[3525] = 16'h732f;
mem_array[3524] = 16'hbd71;
mem_array[3527] = 16'h8650;
mem_array[3526] = 16'hbd80;
mem_array[3529] = 16'hd238;
mem_array[3528] = 16'h3b60;
mem_array[3531] = 16'h583e;
mem_array[3530] = 16'hbcf5;
mem_array[3533] = 16'hc65d;
mem_array[3532] = 16'h3c1b;
mem_array[3535] = 16'hcd16;
mem_array[3534] = 16'h3d0d;
mem_array[3537] = 16'hc752;
mem_array[3536] = 16'h3d43;
mem_array[3539] = 16'h0264;
mem_array[3538] = 16'h3cda;
mem_array[3541] = 16'hc5fa;
mem_array[3540] = 16'hbdc6;
mem_array[3543] = 16'h983e;
mem_array[3542] = 16'h3c16;
mem_array[3545] = 16'h1ff0;
mem_array[3544] = 16'h3b4d;
mem_array[3547] = 16'haee0;
mem_array[3546] = 16'h3ea2;
mem_array[3549] = 16'h3404;
mem_array[3548] = 16'h3d17;
mem_array[3551] = 16'heefc;
mem_array[3550] = 16'hbdb3;
mem_array[3553] = 16'hc02f;
mem_array[3552] = 16'h3d19;
mem_array[3555] = 16'he75d;
mem_array[3554] = 16'h3e76;
mem_array[3557] = 16'h3e6c;
mem_array[3556] = 16'hbc1f;
mem_array[3559] = 16'h843c;
mem_array[3558] = 16'hbcbd;
mem_array[3561] = 16'h19e8;
mem_array[3560] = 16'h3c8f;
mem_array[3563] = 16'h1b75;
mem_array[3562] = 16'h3cf0;
mem_array[3565] = 16'h3f24;
mem_array[3564] = 16'h3ecf;
mem_array[3567] = 16'h4292;
mem_array[3566] = 16'h3d10;
mem_array[3569] = 16'hcb75;
mem_array[3568] = 16'h3cc4;
mem_array[3571] = 16'h51a6;
mem_array[3570] = 16'hbea0;
mem_array[3573] = 16'h47fc;
mem_array[3572] = 16'hbccf;
mem_array[3575] = 16'h5ca1;
mem_array[3574] = 16'hbd89;
mem_array[3577] = 16'hf974;
mem_array[3576] = 16'hbdf9;
mem_array[3579] = 16'h2cfb;
mem_array[3578] = 16'hbeac;
mem_array[3581] = 16'h025c;
mem_array[3580] = 16'h3d86;
mem_array[3583] = 16'h3f71;
mem_array[3582] = 16'h3cdf;
mem_array[3585] = 16'hdb0d;
mem_array[3584] = 16'h3cca;
mem_array[3587] = 16'h3e06;
mem_array[3586] = 16'h3dba;
mem_array[3589] = 16'h7842;
mem_array[3588] = 16'h3a2c;
mem_array[3591] = 16'hbbdf;
mem_array[3590] = 16'h3d8e;
mem_array[3593] = 16'hf604;
mem_array[3592] = 16'h3d2b;
mem_array[3595] = 16'hfd65;
mem_array[3594] = 16'h3bd2;
mem_array[3597] = 16'h1c33;
mem_array[3596] = 16'hbd22;
mem_array[3599] = 16'heacc;
mem_array[3598] = 16'hbecb;
mem_array[3601] = 16'h83b9;
mem_array[3600] = 16'h3c78;
mem_array[3603] = 16'h7cfa;
mem_array[3602] = 16'hbc93;
mem_array[3605] = 16'h7d8b;
mem_array[3604] = 16'hbbd5;
mem_array[3607] = 16'h0736;
mem_array[3606] = 16'h3e89;
mem_array[3609] = 16'h1aa2;
mem_array[3608] = 16'hbd21;
mem_array[3611] = 16'h3c10;
mem_array[3610] = 16'h3dd9;
mem_array[3613] = 16'ha6e5;
mem_array[3612] = 16'h3b95;
mem_array[3615] = 16'h2635;
mem_array[3614] = 16'h3e52;
mem_array[3617] = 16'h9c77;
mem_array[3616] = 16'hbce5;
mem_array[3619] = 16'h4158;
mem_array[3618] = 16'hbd32;
mem_array[3621] = 16'hae16;
mem_array[3620] = 16'hbcef;
mem_array[3623] = 16'hfa5a;
mem_array[3622] = 16'h3cf8;
mem_array[3625] = 16'he96a;
mem_array[3624] = 16'h3eba;
mem_array[3627] = 16'h6965;
mem_array[3626] = 16'hbc37;
mem_array[3629] = 16'h7b3a;
mem_array[3628] = 16'hbc7b;
mem_array[3631] = 16'hf063;
mem_array[3630] = 16'hbeb7;
mem_array[3633] = 16'hbc73;
mem_array[3632] = 16'hbd42;
mem_array[3635] = 16'h35eb;
mem_array[3634] = 16'h3c93;
mem_array[3637] = 16'h251d;
mem_array[3636] = 16'hbded;
mem_array[3639] = 16'h05da;
mem_array[3638] = 16'hbe74;
mem_array[3641] = 16'h7eee;
mem_array[3640] = 16'hbc9e;
mem_array[3643] = 16'h946c;
mem_array[3642] = 16'h3de2;
mem_array[3645] = 16'h6b19;
mem_array[3644] = 16'hbc6a;
mem_array[3647] = 16'h4e8a;
mem_array[3646] = 16'h3bbc;
mem_array[3649] = 16'h5e08;
mem_array[3648] = 16'h3dab;
mem_array[3651] = 16'h7973;
mem_array[3650] = 16'hbd90;
mem_array[3653] = 16'hc6c0;
mem_array[3652] = 16'h3d75;
mem_array[3655] = 16'h06d0;
mem_array[3654] = 16'h3b4f;
mem_array[3657] = 16'hb71c;
mem_array[3656] = 16'hbcab;
mem_array[3659] = 16'hf6cf;
mem_array[3658] = 16'hbeba;
mem_array[3661] = 16'h01e4;
mem_array[3660] = 16'hbce1;
mem_array[3663] = 16'he874;
mem_array[3662] = 16'hbd16;
mem_array[3665] = 16'hc9a1;
mem_array[3664] = 16'h3da4;
mem_array[3667] = 16'h30ab;
mem_array[3666] = 16'hbd8b;
mem_array[3669] = 16'h75c2;
mem_array[3668] = 16'hbd97;
mem_array[3671] = 16'ha77b;
mem_array[3670] = 16'h3d2a;
mem_array[3673] = 16'he78b;
mem_array[3672] = 16'hbd0d;
mem_array[3675] = 16'h5b70;
mem_array[3674] = 16'hbdff;
mem_array[3677] = 16'h7093;
mem_array[3676] = 16'hbdda;
mem_array[3679] = 16'h85da;
mem_array[3678] = 16'h3bd0;
mem_array[3681] = 16'h6388;
mem_array[3680] = 16'hbd5b;
mem_array[3683] = 16'hc58e;
mem_array[3682] = 16'hbd06;
mem_array[3685] = 16'hd14c;
mem_array[3684] = 16'h3e2c;
mem_array[3687] = 16'h42c7;
mem_array[3686] = 16'h3e4b;
mem_array[3689] = 16'h9d54;
mem_array[3688] = 16'h3ddc;
mem_array[3691] = 16'h0067;
mem_array[3690] = 16'hbd42;
mem_array[3693] = 16'hd29c;
mem_array[3692] = 16'h3df1;
mem_array[3695] = 16'hfda7;
mem_array[3694] = 16'hbd28;
mem_array[3697] = 16'h8fce;
mem_array[3696] = 16'hbd75;
mem_array[3699] = 16'h4ba4;
mem_array[3698] = 16'hbe3b;
mem_array[3701] = 16'hf6b1;
mem_array[3700] = 16'h3cc9;
mem_array[3703] = 16'hb567;
mem_array[3702] = 16'h3dc8;
mem_array[3705] = 16'h68f3;
mem_array[3704] = 16'h3d36;
mem_array[3707] = 16'h83bd;
mem_array[3706] = 16'hbd4a;
mem_array[3709] = 16'he983;
mem_array[3708] = 16'h3e06;
mem_array[3711] = 16'h0ec9;
mem_array[3710] = 16'hbdc8;
mem_array[3713] = 16'he6f2;
mem_array[3712] = 16'h3e2c;
mem_array[3715] = 16'h243c;
mem_array[3714] = 16'hbd32;
mem_array[3717] = 16'h0c73;
mem_array[3716] = 16'hbcb3;
mem_array[3719] = 16'he313;
mem_array[3718] = 16'hbe5c;
mem_array[3721] = 16'h9b16;
mem_array[3720] = 16'h3dbf;
mem_array[3723] = 16'h4fb7;
mem_array[3722] = 16'h3ddb;
mem_array[3725] = 16'h7a9e;
mem_array[3724] = 16'h3eb3;
mem_array[3727] = 16'hc278;
mem_array[3726] = 16'hbdf7;
mem_array[3729] = 16'h4b0b;
mem_array[3728] = 16'hbdc6;
mem_array[3731] = 16'hb267;
mem_array[3730] = 16'h3db3;
mem_array[3733] = 16'h5829;
mem_array[3732] = 16'hbd9e;
mem_array[3735] = 16'he8be;
mem_array[3734] = 16'hbde1;
mem_array[3737] = 16'h3fc6;
mem_array[3736] = 16'hbd9c;
mem_array[3739] = 16'h53e4;
mem_array[3738] = 16'hbdc7;
mem_array[3741] = 16'h9800;
mem_array[3740] = 16'hbd43;
mem_array[3743] = 16'h59e3;
mem_array[3742] = 16'hbdc9;
mem_array[3745] = 16'h0351;
mem_array[3744] = 16'h3e9e;
mem_array[3747] = 16'h6923;
mem_array[3746] = 16'h3eb7;
mem_array[3749] = 16'h65c8;
mem_array[3748] = 16'h3e0e;
mem_array[3751] = 16'hf327;
mem_array[3750] = 16'hbe3b;
mem_array[3753] = 16'h748a;
mem_array[3752] = 16'h3e84;
mem_array[3755] = 16'hd792;
mem_array[3754] = 16'hbe30;
mem_array[3757] = 16'h1bb0;
mem_array[3756] = 16'hbe60;
mem_array[3759] = 16'hc0a5;
mem_array[3758] = 16'hbe55;
mem_array[3761] = 16'h50ac;
mem_array[3760] = 16'hbd24;
mem_array[3763] = 16'h2040;
mem_array[3762] = 16'h3ea7;
mem_array[3765] = 16'hac96;
mem_array[3764] = 16'hbdc1;
mem_array[3767] = 16'hb50e;
mem_array[3766] = 16'h3f12;
mem_array[3769] = 16'h0dba;
mem_array[3768] = 16'h3d46;
mem_array[3771] = 16'h8674;
mem_array[3770] = 16'hbd5a;
mem_array[3773] = 16'h7d72;
mem_array[3772] = 16'h3e1a;
mem_array[3775] = 16'h8efc;
mem_array[3774] = 16'hbc89;
mem_array[3777] = 16'h44a1;
mem_array[3776] = 16'hbe37;
mem_array[3779] = 16'h70b8;
mem_array[3778] = 16'hbec9;
mem_array[3781] = 16'ha4ad;
mem_array[3780] = 16'h3d94;
mem_array[3783] = 16'hd517;
mem_array[3782] = 16'h3e03;
mem_array[3785] = 16'h5eb0;
mem_array[3784] = 16'h3e6e;
mem_array[3787] = 16'ha8bd;
mem_array[3786] = 16'hbe94;
mem_array[3789] = 16'hf1f9;
mem_array[3788] = 16'hbe2b;
mem_array[3791] = 16'h8a92;
mem_array[3790] = 16'h3d30;
mem_array[3793] = 16'h4a4b;
mem_array[3792] = 16'h3ef0;
mem_array[3795] = 16'h1e23;
mem_array[3794] = 16'h3f3c;
mem_array[3797] = 16'h03f3;
mem_array[3796] = 16'hbe65;
mem_array[3799] = 16'hb03a;
mem_array[3798] = 16'hbccc;
mem_array[3801] = 16'hc69e;
mem_array[3800] = 16'h3d2e;
mem_array[3803] = 16'h0b57;
mem_array[3802] = 16'hbd0d;
mem_array[3805] = 16'h6afc;
mem_array[3804] = 16'h3e3a;
mem_array[3807] = 16'h2f3a;
mem_array[3806] = 16'h3f73;
mem_array[3809] = 16'hfa29;
mem_array[3808] = 16'h3ea0;
mem_array[3811] = 16'h0838;
mem_array[3810] = 16'hbcd3;
mem_array[3813] = 16'h7424;
mem_array[3812] = 16'h3ed1;
mem_array[3815] = 16'h9f8b;
mem_array[3814] = 16'hbdc2;
mem_array[3817] = 16'h8cdb;
mem_array[3816] = 16'hbe94;
mem_array[3819] = 16'hc8e9;
mem_array[3818] = 16'hbebf;
mem_array[3821] = 16'h5c39;
mem_array[3820] = 16'hbde6;
mem_array[3823] = 16'hd7eb;
mem_array[3822] = 16'h3e98;
mem_array[3825] = 16'h9798;
mem_array[3824] = 16'hbe79;
mem_array[3827] = 16'hca07;
mem_array[3826] = 16'h3f28;
mem_array[3829] = 16'h203d;
mem_array[3828] = 16'h3e01;
mem_array[3831] = 16'hd80c;
mem_array[3830] = 16'hbc87;
mem_array[3833] = 16'h4842;
mem_array[3832] = 16'hba52;
mem_array[3835] = 16'h2eac;
mem_array[3834] = 16'hbd3c;
mem_array[3837] = 16'hb135;
mem_array[3836] = 16'h3e1e;
mem_array[3839] = 16'h0dce;
mem_array[3838] = 16'hbe95;
mem_array[3841] = 16'h6798;
mem_array[3840] = 16'hbce0;
mem_array[3843] = 16'h7477;
mem_array[3842] = 16'h3cfd;
mem_array[3845] = 16'h29cb;
mem_array[3844] = 16'h3e7c;
mem_array[3847] = 16'hb8f1;
mem_array[3846] = 16'h3e7f;
mem_array[3849] = 16'h9a50;
mem_array[3848] = 16'hbf0b;
mem_array[3851] = 16'hea22;
mem_array[3850] = 16'hbf45;
mem_array[3853] = 16'h1fc2;
mem_array[3852] = 16'h3f29;
mem_array[3855] = 16'h2455;
mem_array[3854] = 16'h3eb2;
mem_array[3857] = 16'h2404;
mem_array[3856] = 16'h3e2e;
mem_array[3859] = 16'hcf81;
mem_array[3858] = 16'h3f50;
mem_array[3861] = 16'h6d84;
mem_array[3860] = 16'hbab6;
mem_array[3863] = 16'h9532;
mem_array[3862] = 16'h3dd8;
mem_array[3865] = 16'haba7;
mem_array[3864] = 16'h3f53;
mem_array[3867] = 16'hc341;
mem_array[3866] = 16'h3e09;
mem_array[3869] = 16'h3521;
mem_array[3868] = 16'h3db2;
mem_array[3871] = 16'h83bf;
mem_array[3870] = 16'hbbd6;
mem_array[3873] = 16'hab0b;
mem_array[3872] = 16'h3fe7;
mem_array[3875] = 16'h8c01;
mem_array[3874] = 16'hbe96;
mem_array[3877] = 16'h84d6;
mem_array[3876] = 16'hbe2c;
mem_array[3879] = 16'hd41b;
mem_array[3878] = 16'h3d57;
mem_array[3881] = 16'h02af;
mem_array[3880] = 16'hbe26;
mem_array[3883] = 16'hd3ee;
mem_array[3882] = 16'hbeef;
mem_array[3885] = 16'hf1d7;
mem_array[3884] = 16'hbe88;
mem_array[3887] = 16'hf8de;
mem_array[3886] = 16'h3f42;
mem_array[3889] = 16'h3984;
mem_array[3888] = 16'h3f24;
mem_array[3891] = 16'h0c0d;
mem_array[3890] = 16'hbdc6;
mem_array[3893] = 16'h5d1c;
mem_array[3892] = 16'hbe12;
mem_array[3895] = 16'haf67;
mem_array[3894] = 16'hbe69;
mem_array[3897] = 16'ha806;
mem_array[3896] = 16'h3e9c;
mem_array[3899] = 16'hf019;
mem_array[3898] = 16'hbe37;
mem_array[3901] = 16'ha91f;
mem_array[3900] = 16'hbb19;
mem_array[3903] = 16'hcf29;
mem_array[3902] = 16'hbe09;
mem_array[3905] = 16'h5f6a;
mem_array[3904] = 16'hbd66;
mem_array[3907] = 16'h5931;
mem_array[3906] = 16'hbff2;
mem_array[3909] = 16'hc646;
mem_array[3908] = 16'h3ec4;
mem_array[3911] = 16'ha0e2;
mem_array[3910] = 16'hbf15;
mem_array[3913] = 16'h51e7;
mem_array[3912] = 16'h3f38;
mem_array[3915] = 16'h0975;
mem_array[3914] = 16'hbe35;
mem_array[3917] = 16'h40a8;
mem_array[3916] = 16'h3ef2;
mem_array[3919] = 16'h9e9e;
mem_array[3918] = 16'h3e94;
mem_array[3921] = 16'h4798;
mem_array[3920] = 16'hbd11;
mem_array[3923] = 16'ha2cb;
mem_array[3922] = 16'h3d6f;
mem_array[3925] = 16'h2dd3;
mem_array[3924] = 16'h3f9f;
mem_array[3927] = 16'h4e88;
mem_array[3926] = 16'h3ece;
mem_array[3929] = 16'h2f0a;
mem_array[3928] = 16'h3edf;
mem_array[3931] = 16'hb839;
mem_array[3930] = 16'hbf01;
mem_array[3933] = 16'h2286;
mem_array[3932] = 16'h3fd2;
mem_array[3935] = 16'hfae6;
mem_array[3934] = 16'hbe87;
mem_array[3937] = 16'h5b6e;
mem_array[3936] = 16'hbe80;
mem_array[3939] = 16'h3d95;
mem_array[3938] = 16'h3ec3;
mem_array[3941] = 16'hb57b;
mem_array[3940] = 16'hbe18;
mem_array[3943] = 16'hf407;
mem_array[3942] = 16'hbf0c;
mem_array[3945] = 16'hf07e;
mem_array[3944] = 16'hbf27;
mem_array[3947] = 16'h8f9d;
mem_array[3946] = 16'h3fee;
mem_array[3949] = 16'h12ef;
mem_array[3948] = 16'h3e45;
mem_array[3951] = 16'h4f0f;
mem_array[3950] = 16'hbb80;
mem_array[3953] = 16'h0cae;
mem_array[3952] = 16'hbf10;
mem_array[3955] = 16'h8f72;
mem_array[3954] = 16'hbeba;
mem_array[3957] = 16'h8261;
mem_array[3956] = 16'h3f6b;
mem_array[3959] = 16'h7f6d;
mem_array[3958] = 16'h3e6e;
mem_array[3961] = 16'h5468;
mem_array[3960] = 16'h3db7;
mem_array[3963] = 16'h5dc2;
mem_array[3962] = 16'hbe23;
mem_array[3965] = 16'h9fb5;
mem_array[3964] = 16'h3e64;
mem_array[3967] = 16'h2c89;
mem_array[3966] = 16'hbe40;
mem_array[3969] = 16'he109;
mem_array[3968] = 16'hbf0d;
mem_array[3971] = 16'hde25;
mem_array[3970] = 16'hbf7c;
mem_array[3973] = 16'hc1fc;
mem_array[3972] = 16'h3e3d;
mem_array[3975] = 16'hf7e4;
mem_array[3974] = 16'h3f83;
mem_array[3977] = 16'h9c3a;
mem_array[3976] = 16'h3d3d;
mem_array[3979] = 16'hea74;
mem_array[3978] = 16'h3f0c;
mem_array[3981] = 16'h674f;
mem_array[3980] = 16'hbdcc;
mem_array[3983] = 16'h40e9;
mem_array[3982] = 16'h3c7a;
mem_array[3985] = 16'h487d;
mem_array[3984] = 16'h3f99;
mem_array[3987] = 16'hedae;
mem_array[3986] = 16'hbbf8;
mem_array[3989] = 16'h86eb;
mem_array[3988] = 16'h3f3f;
mem_array[3991] = 16'h76dd;
mem_array[3990] = 16'hbf22;
mem_array[3993] = 16'h4198;
mem_array[3992] = 16'h3f37;
mem_array[3995] = 16'hb05b;
mem_array[3994] = 16'hbf06;
mem_array[3997] = 16'h09c3;
mem_array[3996] = 16'hbf30;
mem_array[3999] = 16'hbc64;
mem_array[3998] = 16'h3e78;
mem_array[4001] = 16'hd049;
mem_array[4000] = 16'hbf5c;
mem_array[4003] = 16'h82ff;
mem_array[4002] = 16'h3db7;
mem_array[4005] = 16'h2263;
mem_array[4004] = 16'hbea2;
mem_array[4007] = 16'h0e98;
mem_array[4006] = 16'h3fd3;
mem_array[4009] = 16'ha27c;
mem_array[4008] = 16'h3f12;
mem_array[4011] = 16'h8aee;
mem_array[4010] = 16'hbd16;
mem_array[4013] = 16'h5564;
mem_array[4012] = 16'hbe6a;
mem_array[4015] = 16'h4031;
mem_array[4014] = 16'hbe92;
mem_array[4017] = 16'h54ff;
mem_array[4016] = 16'h3f81;
mem_array[4019] = 16'h652e;
mem_array[4018] = 16'h3ed7;
mem_array[4021] = 16'h22c6;
mem_array[4020] = 16'hbc91;
mem_array[4023] = 16'h11dd;
mem_array[4022] = 16'hbeb3;
mem_array[4025] = 16'hb8d1;
mem_array[4024] = 16'h3f29;
mem_array[4027] = 16'he24c;
mem_array[4026] = 16'hbf62;
mem_array[4029] = 16'h3fef;
mem_array[4028] = 16'hbe3f;
mem_array[4031] = 16'h0079;
mem_array[4030] = 16'hbf0f;
mem_array[4033] = 16'hfdc3;
mem_array[4032] = 16'h3f5e;
mem_array[4035] = 16'h66e2;
mem_array[4034] = 16'h3f6b;
mem_array[4037] = 16'heb10;
mem_array[4036] = 16'hbd90;
mem_array[4039] = 16'ha6d8;
mem_array[4038] = 16'h3f64;
mem_array[4041] = 16'h8d92;
mem_array[4040] = 16'hbd75;
mem_array[4043] = 16'h9329;
mem_array[4042] = 16'hbd87;
mem_array[4045] = 16'ha6de;
mem_array[4044] = 16'h3f6f;
mem_array[4047] = 16'h0b7a;
mem_array[4046] = 16'hbd94;
mem_array[4049] = 16'h7234;
mem_array[4048] = 16'hbd32;
mem_array[4051] = 16'hd851;
mem_array[4050] = 16'hbf54;
mem_array[4053] = 16'he68b;
mem_array[4052] = 16'h3dbc;
mem_array[4055] = 16'h53b3;
mem_array[4054] = 16'hbfbe;
mem_array[4057] = 16'h76a4;
mem_array[4056] = 16'hbfcc;
mem_array[4059] = 16'h1845;
mem_array[4058] = 16'h3e1e;
mem_array[4061] = 16'he105;
mem_array[4060] = 16'hbf69;
mem_array[4063] = 16'h8ad8;
mem_array[4062] = 16'hbd4f;
mem_array[4065] = 16'hf763;
mem_array[4064] = 16'h3e03;
mem_array[4067] = 16'hbc12;
mem_array[4066] = 16'h3fd0;
mem_array[4069] = 16'h80ab;
mem_array[4068] = 16'h3eca;
mem_array[4071] = 16'hca95;
mem_array[4070] = 16'hbe00;
mem_array[4073] = 16'hc731;
mem_array[4072] = 16'h3e85;
mem_array[4075] = 16'h9db0;
mem_array[4074] = 16'hbf13;
mem_array[4077] = 16'h6c50;
mem_array[4076] = 16'h3f91;
mem_array[4079] = 16'h67dd;
mem_array[4078] = 16'h3f3e;
mem_array[4081] = 16'h797a;
mem_array[4080] = 16'hbed0;
mem_array[4083] = 16'he032;
mem_array[4082] = 16'hbe2d;
mem_array[4085] = 16'h2ab8;
mem_array[4084] = 16'h3fc4;
mem_array[4087] = 16'h6b15;
mem_array[4086] = 16'h3cc5;
mem_array[4089] = 16'h72d3;
mem_array[4088] = 16'hbd5b;
mem_array[4091] = 16'hbad6;
mem_array[4090] = 16'hbfcf;
mem_array[4093] = 16'h5bc6;
mem_array[4092] = 16'h3e87;
mem_array[4095] = 16'he7b5;
mem_array[4094] = 16'h3d67;
mem_array[4097] = 16'h4635;
mem_array[4096] = 16'hbdff;
mem_array[4099] = 16'h5f36;
mem_array[4098] = 16'h3e2a;
mem_array[4101] = 16'h654d;
mem_array[4100] = 16'hbdb2;
mem_array[4103] = 16'hbf0d;
mem_array[4102] = 16'hbd3a;
mem_array[4105] = 16'h4c3f;
mem_array[4104] = 16'h3fe6;
mem_array[4107] = 16'h27fa;
mem_array[4106] = 16'hbe5a;
mem_array[4109] = 16'hdf96;
mem_array[4108] = 16'h3d34;
mem_array[4111] = 16'h607c;
mem_array[4110] = 16'h3eca;
mem_array[4113] = 16'hc030;
mem_array[4112] = 16'h3eac;
mem_array[4115] = 16'h13ab;
mem_array[4114] = 16'hbf8a;
mem_array[4117] = 16'h6f9f;
mem_array[4116] = 16'hbfd8;
mem_array[4119] = 16'h05d9;
mem_array[4118] = 16'hbf09;
mem_array[4121] = 16'hb10b;
mem_array[4120] = 16'hbf10;
mem_array[4123] = 16'hd6b3;
mem_array[4122] = 16'h3ec6;
mem_array[4125] = 16'hd526;
mem_array[4124] = 16'hbfc3;
mem_array[4127] = 16'h8ee6;
mem_array[4126] = 16'h402a;
mem_array[4129] = 16'h661a;
mem_array[4128] = 16'hbece;
mem_array[4131] = 16'h6f7d;
mem_array[4130] = 16'hbd94;
mem_array[4133] = 16'h993c;
mem_array[4132] = 16'h3f77;
mem_array[4135] = 16'h743d;
mem_array[4134] = 16'hbe58;
mem_array[4137] = 16'h8954;
mem_array[4136] = 16'hbdd0;
mem_array[4139] = 16'hce87;
mem_array[4138] = 16'h3efe;
mem_array[4141] = 16'h6fa1;
mem_array[4140] = 16'hbec5;
mem_array[4143] = 16'hed17;
mem_array[4142] = 16'hbeb9;
mem_array[4145] = 16'h121f;
mem_array[4144] = 16'h3ea3;
mem_array[4147] = 16'h15e9;
mem_array[4146] = 16'hbee6;
mem_array[4149] = 16'ha576;
mem_array[4148] = 16'hbe84;
mem_array[4151] = 16'hf80f;
mem_array[4150] = 16'h3e1c;
mem_array[4153] = 16'ha461;
mem_array[4152] = 16'h3e6b;
mem_array[4155] = 16'h1132;
mem_array[4154] = 16'hbc83;
mem_array[4157] = 16'h45b5;
mem_array[4156] = 16'h3db2;
mem_array[4159] = 16'h7538;
mem_array[4158] = 16'h3f62;
mem_array[4161] = 16'h2e56;
mem_array[4160] = 16'h3d9b;
mem_array[4163] = 16'h5e3f;
mem_array[4162] = 16'hbdcb;
mem_array[4165] = 16'h3f15;
mem_array[4164] = 16'h3f7b;
mem_array[4167] = 16'hd768;
mem_array[4166] = 16'h3ea5;
mem_array[4169] = 16'h0b76;
mem_array[4168] = 16'h3ea1;
mem_array[4171] = 16'hec7a;
mem_array[4170] = 16'hbe83;
mem_array[4173] = 16'hb71b;
mem_array[4172] = 16'h3f95;
mem_array[4175] = 16'hcd27;
mem_array[4174] = 16'hbf82;
mem_array[4177] = 16'he681;
mem_array[4176] = 16'hbfd5;
mem_array[4179] = 16'hcb49;
mem_array[4178] = 16'hbf05;
mem_array[4181] = 16'haa0a;
mem_array[4180] = 16'hbf1f;
mem_array[4183] = 16'hdd64;
mem_array[4182] = 16'h3b25;
mem_array[4185] = 16'h4bb7;
mem_array[4184] = 16'hbfb0;
mem_array[4187] = 16'h5f61;
mem_array[4186] = 16'h4002;
mem_array[4189] = 16'had4b;
mem_array[4188] = 16'h3f01;
mem_array[4191] = 16'h529a;
mem_array[4190] = 16'hbcfc;
mem_array[4193] = 16'h16ed;
mem_array[4192] = 16'h3d52;
mem_array[4195] = 16'ha826;
mem_array[4194] = 16'h3b1d;
mem_array[4197] = 16'hc824;
mem_array[4196] = 16'h3f80;
mem_array[4199] = 16'hec2b;
mem_array[4198] = 16'h3f07;
mem_array[4201] = 16'h1a17;
mem_array[4200] = 16'hbef7;
mem_array[4203] = 16'h8d79;
mem_array[4202] = 16'hbf4b;
mem_array[4205] = 16'h6e2a;
mem_array[4204] = 16'hbf26;
mem_array[4207] = 16'hcb8b;
mem_array[4206] = 16'hbfb4;
mem_array[4209] = 16'hef7e;
mem_array[4208] = 16'hbead;
mem_array[4211] = 16'h6c45;
mem_array[4210] = 16'h3d9a;
mem_array[4213] = 16'h03cc;
mem_array[4212] = 16'hbf1a;
mem_array[4215] = 16'h9b5d;
mem_array[4214] = 16'h3e26;
mem_array[4217] = 16'h31b5;
mem_array[4216] = 16'hbf38;
mem_array[4219] = 16'h82f1;
mem_array[4218] = 16'h3eb4;
mem_array[4221] = 16'h93e0;
mem_array[4220] = 16'hbd88;
mem_array[4223] = 16'he164;
mem_array[4222] = 16'hbd05;
mem_array[4225] = 16'hfbb5;
mem_array[4224] = 16'h3f07;
mem_array[4227] = 16'hfce4;
mem_array[4226] = 16'hbeb8;
mem_array[4229] = 16'h20a0;
mem_array[4228] = 16'h3f39;
mem_array[4231] = 16'h6ae1;
mem_array[4230] = 16'h3e06;
mem_array[4233] = 16'h5c56;
mem_array[4232] = 16'h3e41;
mem_array[4235] = 16'h149c;
mem_array[4234] = 16'hbfa1;
mem_array[4237] = 16'h864a;
mem_array[4236] = 16'hbfd8;
mem_array[4239] = 16'ha696;
mem_array[4238] = 16'h3f5f;
mem_array[4241] = 16'h97bc;
mem_array[4240] = 16'hbf98;
mem_array[4243] = 16'h8484;
mem_array[4242] = 16'hbe52;
mem_array[4245] = 16'h17ff;
mem_array[4244] = 16'hbde6;
mem_array[4247] = 16'h5fe5;
mem_array[4246] = 16'h3f91;
mem_array[4249] = 16'hde29;
mem_array[4248] = 16'h3f18;
mem_array[4251] = 16'h1a00;
mem_array[4250] = 16'hbf02;
mem_array[4253] = 16'hcda4;
mem_array[4252] = 16'hbe69;
mem_array[4255] = 16'hd308;
mem_array[4254] = 16'hbeb9;
mem_array[4257] = 16'h34a0;
mem_array[4256] = 16'h3f0d;
mem_array[4259] = 16'hafe1;
mem_array[4258] = 16'h3f2b;
mem_array[4261] = 16'h4d45;
mem_array[4260] = 16'hbfc4;
mem_array[4263] = 16'h7f76;
mem_array[4262] = 16'hbf0c;
mem_array[4265] = 16'h8331;
mem_array[4264] = 16'hbf80;
mem_array[4267] = 16'hf3c8;
mem_array[4266] = 16'hbfb5;
mem_array[4269] = 16'hfe9e;
mem_array[4268] = 16'hbe0a;
mem_array[4271] = 16'hc293;
mem_array[4270] = 16'h3ed3;
mem_array[4273] = 16'h9877;
mem_array[4272] = 16'hbf71;
mem_array[4275] = 16'hc5f2;
mem_array[4274] = 16'h3e97;
mem_array[4277] = 16'hb2a8;
mem_array[4276] = 16'hbf17;
mem_array[4279] = 16'hecee;
mem_array[4278] = 16'h3ea5;
mem_array[4281] = 16'he533;
mem_array[4280] = 16'hbd2a;
mem_array[4283] = 16'ha91f;
mem_array[4282] = 16'hbd89;
mem_array[4285] = 16'h6301;
mem_array[4284] = 16'hbf21;
mem_array[4287] = 16'h059e;
mem_array[4286] = 16'hbf7a;
mem_array[4289] = 16'hbc4e;
mem_array[4288] = 16'h3f58;
mem_array[4291] = 16'h576e;
mem_array[4290] = 16'h3f74;
mem_array[4293] = 16'h28e1;
mem_array[4292] = 16'h3ebd;
mem_array[4295] = 16'h5921;
mem_array[4294] = 16'hbf2f;
mem_array[4297] = 16'h31db;
mem_array[4296] = 16'hbf84;
mem_array[4299] = 16'h06ff;
mem_array[4298] = 16'hbd6d;
mem_array[4301] = 16'hc825;
mem_array[4300] = 16'hbeaf;
mem_array[4303] = 16'hb029;
mem_array[4302] = 16'hbe1c;
mem_array[4305] = 16'h1e1d;
mem_array[4304] = 16'h3dbb;
mem_array[4307] = 16'h0ff1;
mem_array[4306] = 16'h3f18;
mem_array[4309] = 16'h78fb;
mem_array[4308] = 16'h3ee4;
mem_array[4311] = 16'h39cf;
mem_array[4310] = 16'hbf59;
mem_array[4313] = 16'h35ae;
mem_array[4312] = 16'h3df3;
mem_array[4315] = 16'h5327;
mem_array[4314] = 16'h3dd8;
mem_array[4317] = 16'h6572;
mem_array[4316] = 16'h3f2a;
mem_array[4319] = 16'h6341;
mem_array[4318] = 16'h3e73;
mem_array[4321] = 16'h1572;
mem_array[4320] = 16'hbffa;
mem_array[4323] = 16'hc308;
mem_array[4322] = 16'hbf2c;
mem_array[4325] = 16'hcc0c;
mem_array[4324] = 16'hbfa0;
mem_array[4327] = 16'h44f2;
mem_array[4326] = 16'hbfc2;
mem_array[4329] = 16'hbf3a;
mem_array[4328] = 16'hbe47;
mem_array[4331] = 16'h651c;
mem_array[4330] = 16'h3e67;
mem_array[4333] = 16'h085f;
mem_array[4332] = 16'hbf73;
mem_array[4335] = 16'h54e7;
mem_array[4334] = 16'h3e92;
mem_array[4337] = 16'h457a;
mem_array[4336] = 16'h3e87;
mem_array[4339] = 16'he245;
mem_array[4338] = 16'h3f76;
mem_array[4341] = 16'h1489;
mem_array[4340] = 16'hbd89;
mem_array[4343] = 16'h3fea;
mem_array[4342] = 16'hbc11;
mem_array[4345] = 16'h79c9;
mem_array[4344] = 16'hbd41;
mem_array[4347] = 16'h83b9;
mem_array[4346] = 16'hbf2d;
mem_array[4349] = 16'h8926;
mem_array[4348] = 16'h3e91;
mem_array[4351] = 16'h3201;
mem_array[4350] = 16'h3ec4;
mem_array[4353] = 16'h4252;
mem_array[4352] = 16'hbd9c;
mem_array[4355] = 16'hf815;
mem_array[4354] = 16'hbd23;
mem_array[4357] = 16'haacd;
mem_array[4356] = 16'hbfce;
mem_array[4359] = 16'hd741;
mem_array[4358] = 16'h3cee;
mem_array[4361] = 16'h9848;
mem_array[4360] = 16'hbe90;
mem_array[4363] = 16'h6d99;
mem_array[4362] = 16'h3e30;
mem_array[4365] = 16'he61a;
mem_array[4364] = 16'h3ea3;
mem_array[4367] = 16'h6dd8;
mem_array[4366] = 16'h3e42;
mem_array[4369] = 16'hcfc4;
mem_array[4368] = 16'hbeb2;
mem_array[4371] = 16'hc5fe;
mem_array[4370] = 16'hbf14;
mem_array[4373] = 16'h8fe8;
mem_array[4372] = 16'hbebb;
mem_array[4375] = 16'h4995;
mem_array[4374] = 16'h3d80;
mem_array[4377] = 16'h15df;
mem_array[4376] = 16'h3f67;
mem_array[4379] = 16'had61;
mem_array[4378] = 16'h3e33;
mem_array[4381] = 16'h6023;
mem_array[4380] = 16'hbfd3;
mem_array[4383] = 16'h2903;
mem_array[4382] = 16'hbf2f;
mem_array[4385] = 16'hbe1e;
mem_array[4384] = 16'hbfb9;
mem_array[4387] = 16'hc9e3;
mem_array[4386] = 16'hbf72;
mem_array[4389] = 16'ha3ef;
mem_array[4388] = 16'hbf1b;
mem_array[4391] = 16'h246a;
mem_array[4390] = 16'hbedf;
mem_array[4393] = 16'hce87;
mem_array[4392] = 16'hbf78;
mem_array[4395] = 16'h6bce;
mem_array[4394] = 16'hbeb8;
mem_array[4397] = 16'h5292;
mem_array[4396] = 16'hbe6c;
mem_array[4399] = 16'h4489;
mem_array[4398] = 16'hbf90;
mem_array[4401] = 16'he2a2;
mem_array[4400] = 16'hbe0b;
mem_array[4403] = 16'h5d5a;
mem_array[4402] = 16'h3d3d;
mem_array[4405] = 16'heffa;
mem_array[4404] = 16'hbb22;
mem_array[4407] = 16'h4c09;
mem_array[4406] = 16'hbef5;
mem_array[4409] = 16'h6fd8;
mem_array[4408] = 16'h3d7e;
mem_array[4411] = 16'h9d93;
mem_array[4410] = 16'hbeb5;
mem_array[4413] = 16'h6afe;
mem_array[4412] = 16'hbed7;
mem_array[4415] = 16'h4ff0;
mem_array[4414] = 16'hbeb4;
mem_array[4417] = 16'he435;
mem_array[4416] = 16'hbf8c;
mem_array[4419] = 16'hc56f;
mem_array[4418] = 16'h3e1e;
mem_array[4421] = 16'h119c;
mem_array[4420] = 16'hbf86;
mem_array[4423] = 16'h5d74;
mem_array[4422] = 16'h3ec7;
mem_array[4425] = 16'h368c;
mem_array[4424] = 16'h3edc;
mem_array[4427] = 16'h47a6;
mem_array[4426] = 16'h3f7d;
mem_array[4429] = 16'h8a3b;
mem_array[4428] = 16'hbeb2;
mem_array[4431] = 16'h9b2e;
mem_array[4430] = 16'hbefc;
mem_array[4433] = 16'h97fc;
mem_array[4432] = 16'hbf31;
mem_array[4435] = 16'h6662;
mem_array[4434] = 16'h3f29;
mem_array[4437] = 16'h2e54;
mem_array[4436] = 16'h3f06;
mem_array[4439] = 16'h55a4;
mem_array[4438] = 16'hbe2d;
mem_array[4441] = 16'h5ea9;
mem_array[4440] = 16'hbfc0;
mem_array[4443] = 16'h578b;
mem_array[4442] = 16'hbebd;
mem_array[4445] = 16'h028d;
mem_array[4444] = 16'hbf96;
mem_array[4447] = 16'hddab;
mem_array[4446] = 16'hbfd1;
mem_array[4449] = 16'h3de7;
mem_array[4448] = 16'hbf28;
mem_array[4451] = 16'h6fd1;
mem_array[4450] = 16'h3ef7;
mem_array[4453] = 16'h5fd3;
mem_array[4452] = 16'hbff1;
mem_array[4455] = 16'h382f;
mem_array[4454] = 16'h3e33;
mem_array[4457] = 16'h0b2a;
mem_array[4456] = 16'h3cb1;
mem_array[4459] = 16'h785a;
mem_array[4458] = 16'hbfe5;
mem_array[4461] = 16'h21e3;
mem_array[4460] = 16'h3d24;
mem_array[4463] = 16'h714f;
mem_array[4462] = 16'hbd4e;
mem_array[4465] = 16'h1e4c;
mem_array[4464] = 16'hbe5b;
mem_array[4467] = 16'h159a;
mem_array[4466] = 16'hbf54;
mem_array[4469] = 16'h311c;
mem_array[4468] = 16'hbe01;
mem_array[4471] = 16'h5ad7;
mem_array[4470] = 16'hbf0a;
mem_array[4473] = 16'h693b;
mem_array[4472] = 16'hbfd2;
mem_array[4475] = 16'h83ec;
mem_array[4474] = 16'hbf37;
mem_array[4477] = 16'h3623;
mem_array[4476] = 16'hbfa4;
mem_array[4479] = 16'hacfd;
mem_array[4478] = 16'hbf3c;
mem_array[4481] = 16'h3253;
mem_array[4480] = 16'hbf7d;
mem_array[4483] = 16'h4b1b;
mem_array[4482] = 16'h3f17;
mem_array[4485] = 16'h3da2;
mem_array[4484] = 16'h3e74;
mem_array[4487] = 16'h4773;
mem_array[4486] = 16'h3f5b;
mem_array[4489] = 16'he2fe;
mem_array[4488] = 16'hbeaa;
mem_array[4491] = 16'hc42b;
mem_array[4490] = 16'hbdac;
mem_array[4493] = 16'ha486;
mem_array[4492] = 16'hbe90;
mem_array[4495] = 16'h0036;
mem_array[4494] = 16'h3f9b;
mem_array[4497] = 16'hfc68;
mem_array[4496] = 16'h3e6d;
mem_array[4499] = 16'h137b;
mem_array[4498] = 16'hbf18;
mem_array[4501] = 16'h1fbf;
mem_array[4500] = 16'h3d09;
mem_array[4503] = 16'hfe76;
mem_array[4502] = 16'hbdc1;
mem_array[4505] = 16'h197f;
mem_array[4504] = 16'hbeaa;
mem_array[4507] = 16'h5b0d;
mem_array[4506] = 16'hbff7;
mem_array[4509] = 16'hbf95;
mem_array[4508] = 16'hbee1;
mem_array[4511] = 16'h2b5a;
mem_array[4510] = 16'h3ecb;
mem_array[4513] = 16'hffbc;
mem_array[4512] = 16'hbf98;
mem_array[4515] = 16'hbbed;
mem_array[4514] = 16'hbf27;
mem_array[4517] = 16'he9dc;
mem_array[4516] = 16'hbe19;
mem_array[4519] = 16'h6043;
mem_array[4518] = 16'hbf5f;
mem_array[4521] = 16'he4ce;
mem_array[4520] = 16'h3d22;
mem_array[4523] = 16'h2c48;
mem_array[4522] = 16'hbd41;
mem_array[4525] = 16'he763;
mem_array[4524] = 16'h3efe;
mem_array[4527] = 16'h2836;
mem_array[4526] = 16'hbf9b;
mem_array[4529] = 16'hb6c1;
mem_array[4528] = 16'hbd75;
mem_array[4531] = 16'h5461;
mem_array[4530] = 16'hbf65;
mem_array[4533] = 16'h0f7b;
mem_array[4532] = 16'hbfd3;
mem_array[4535] = 16'h0f9b;
mem_array[4534] = 16'hbed3;
mem_array[4537] = 16'hf794;
mem_array[4536] = 16'hbf9f;
mem_array[4539] = 16'h10c2;
mem_array[4538] = 16'hbe68;
mem_array[4541] = 16'h4ca5;
mem_array[4540] = 16'hbf92;
mem_array[4543] = 16'h6906;
mem_array[4542] = 16'h3f0a;
mem_array[4545] = 16'h544d;
mem_array[4544] = 16'h3f73;
mem_array[4547] = 16'h488e;
mem_array[4546] = 16'h3f90;
mem_array[4549] = 16'h9ecf;
mem_array[4548] = 16'hbee1;
mem_array[4551] = 16'h00bd;
mem_array[4550] = 16'h3d37;
mem_array[4553] = 16'h1774;
mem_array[4552] = 16'hbf08;
mem_array[4555] = 16'h3746;
mem_array[4554] = 16'h3f45;
mem_array[4557] = 16'hccc2;
mem_array[4556] = 16'hbe92;
mem_array[4559] = 16'hed3b;
mem_array[4558] = 16'hbf29;
mem_array[4561] = 16'hff9a;
mem_array[4560] = 16'h3e91;
mem_array[4563] = 16'hda38;
mem_array[4562] = 16'hbd39;
mem_array[4565] = 16'h2c01;
mem_array[4564] = 16'hbf31;
mem_array[4567] = 16'h7dc4;
mem_array[4566] = 16'hbee2;
mem_array[4569] = 16'hca87;
mem_array[4568] = 16'hbeb3;
mem_array[4571] = 16'h4465;
mem_array[4570] = 16'h3e87;
mem_array[4573] = 16'hbcef;
mem_array[4572] = 16'hbf00;
mem_array[4575] = 16'h1ff9;
mem_array[4574] = 16'hbeae;
mem_array[4577] = 16'h1a94;
mem_array[4576] = 16'h3f2e;
mem_array[4579] = 16'h5fb7;
mem_array[4578] = 16'h3de6;
mem_array[4581] = 16'hded2;
mem_array[4580] = 16'h3c36;
mem_array[4583] = 16'h1ee7;
mem_array[4582] = 16'hbdf4;
mem_array[4585] = 16'h0b9f;
mem_array[4584] = 16'hbe49;
mem_array[4587] = 16'h428b;
mem_array[4586] = 16'hbf31;
mem_array[4589] = 16'h23a7;
mem_array[4588] = 16'hbdc3;
mem_array[4591] = 16'had0f;
mem_array[4590] = 16'hbe7e;
mem_array[4593] = 16'h3b81;
mem_array[4592] = 16'hbfe5;
mem_array[4595] = 16'h4789;
mem_array[4594] = 16'hbbc4;
mem_array[4597] = 16'h9979;
mem_array[4596] = 16'hbfa5;
mem_array[4599] = 16'h7e1c;
mem_array[4598] = 16'h3dde;
mem_array[4601] = 16'h06de;
mem_array[4600] = 16'h3f0f;
mem_array[4603] = 16'h831e;
mem_array[4602] = 16'h3f13;
mem_array[4605] = 16'hd8ee;
mem_array[4604] = 16'hbd82;
mem_array[4607] = 16'hfd4c;
mem_array[4606] = 16'h3f21;
mem_array[4609] = 16'h1c71;
mem_array[4608] = 16'h3ed3;
mem_array[4611] = 16'h2ba1;
mem_array[4610] = 16'h3d00;
mem_array[4613] = 16'h619f;
mem_array[4612] = 16'hbd8a;
mem_array[4615] = 16'h0d47;
mem_array[4614] = 16'h3ef6;
mem_array[4617] = 16'h8d6e;
mem_array[4616] = 16'hbe86;
mem_array[4619] = 16'hcdde;
mem_array[4618] = 16'hbe7c;
mem_array[4621] = 16'h731d;
mem_array[4620] = 16'h3e36;
mem_array[4623] = 16'h6e5d;
mem_array[4622] = 16'hbcf4;
mem_array[4625] = 16'hd89f;
mem_array[4624] = 16'hbe58;
mem_array[4627] = 16'h3ff4;
mem_array[4626] = 16'h3e5e;
mem_array[4629] = 16'hf87f;
mem_array[4628] = 16'hbe8f;
mem_array[4631] = 16'h67b5;
mem_array[4630] = 16'hbe24;
mem_array[4633] = 16'h875c;
mem_array[4632] = 16'h3e85;
mem_array[4635] = 16'hcf30;
mem_array[4634] = 16'h3d20;
mem_array[4637] = 16'hfe2a;
mem_array[4636] = 16'h3f17;
mem_array[4639] = 16'hfa5a;
mem_array[4638] = 16'h3e03;
mem_array[4641] = 16'hbc63;
mem_array[4640] = 16'hbd63;
mem_array[4643] = 16'h5926;
mem_array[4642] = 16'h3dc7;
mem_array[4645] = 16'h88f1;
mem_array[4644] = 16'h3dad;
mem_array[4647] = 16'hd088;
mem_array[4646] = 16'h3f8d;
mem_array[4649] = 16'h8b3a;
mem_array[4648] = 16'h3f0f;
mem_array[4651] = 16'h7133;
mem_array[4650] = 16'hbf6e;
mem_array[4653] = 16'h6351;
mem_array[4652] = 16'h3f5e;
mem_array[4655] = 16'hf982;
mem_array[4654] = 16'h3ec5;
mem_array[4657] = 16'h38fe;
mem_array[4656] = 16'hbf1f;
mem_array[4659] = 16'h45ed;
mem_array[4658] = 16'h3e22;
mem_array[4661] = 16'hae89;
mem_array[4660] = 16'h3f37;
mem_array[4663] = 16'hdc6e;
mem_array[4662] = 16'hbe32;
mem_array[4665] = 16'h3321;
mem_array[4664] = 16'h3e5e;
mem_array[4667] = 16'h6d77;
mem_array[4666] = 16'h3ea1;
mem_array[4669] = 16'h651b;
mem_array[4668] = 16'h3f0f;
mem_array[4671] = 16'heb31;
mem_array[4670] = 16'h3c76;
mem_array[4673] = 16'hd81e;
mem_array[4672] = 16'hbca5;
mem_array[4675] = 16'hc3c6;
mem_array[4674] = 16'h3ec8;
mem_array[4677] = 16'h03bd;
mem_array[4676] = 16'h3e5a;
mem_array[4679] = 16'h0398;
mem_array[4678] = 16'hbe3d;
mem_array[4681] = 16'h415e;
mem_array[4680] = 16'h3db6;
mem_array[4683] = 16'he492;
mem_array[4682] = 16'hbba4;
mem_array[4685] = 16'h4efb;
mem_array[4684] = 16'hbda6;
mem_array[4687] = 16'h0188;
mem_array[4686] = 16'h3e3a;
mem_array[4689] = 16'hfef9;
mem_array[4688] = 16'hbe7b;
mem_array[4691] = 16'h90e6;
mem_array[4690] = 16'h3eab;
mem_array[4693] = 16'he6dc;
mem_array[4692] = 16'h3e6d;
mem_array[4695] = 16'ha26b;
mem_array[4694] = 16'h3e92;
mem_array[4697] = 16'h704f;
mem_array[4696] = 16'hbdc3;
mem_array[4699] = 16'hf841;
mem_array[4698] = 16'h3eeb;
mem_array[4701] = 16'h3498;
mem_array[4700] = 16'h3d11;
mem_array[4703] = 16'h367b;
mem_array[4702] = 16'hbc26;
mem_array[4705] = 16'hda2a;
mem_array[4704] = 16'h3e1b;
mem_array[4707] = 16'h8221;
mem_array[4706] = 16'h3d39;
mem_array[4709] = 16'hc698;
mem_array[4708] = 16'h3d1c;
mem_array[4711] = 16'h3df5;
mem_array[4710] = 16'hbf27;
mem_array[4713] = 16'h081a;
mem_array[4712] = 16'hbd74;
mem_array[4715] = 16'h75ab;
mem_array[4714] = 16'h3f2e;
mem_array[4717] = 16'hc389;
mem_array[4716] = 16'hbdb2;
mem_array[4719] = 16'h2672;
mem_array[4718] = 16'h3eaa;
mem_array[4721] = 16'h385e;
mem_array[4720] = 16'h3e46;
mem_array[4723] = 16'h4f37;
mem_array[4722] = 16'hbd80;
mem_array[4725] = 16'hb1c7;
mem_array[4724] = 16'h3dd9;
mem_array[4727] = 16'h28fe;
mem_array[4726] = 16'h3f1b;
mem_array[4729] = 16'h3cfb;
mem_array[4728] = 16'h3e05;
mem_array[4731] = 16'h46f2;
mem_array[4730] = 16'h3c99;
mem_array[4733] = 16'ha68c;
mem_array[4732] = 16'hbecf;
mem_array[4735] = 16'h9092;
mem_array[4734] = 16'h3ea1;
mem_array[4737] = 16'hc310;
mem_array[4736] = 16'hbdb3;
mem_array[4739] = 16'h583a;
mem_array[4738] = 16'h3e96;
mem_array[4741] = 16'h132e;
mem_array[4740] = 16'h3c6e;
mem_array[4743] = 16'h17ef;
mem_array[4742] = 16'h3b4d;
mem_array[4745] = 16'h2986;
mem_array[4744] = 16'h3f7e;
mem_array[4747] = 16'h895b;
mem_array[4746] = 16'h3d86;
mem_array[4749] = 16'h1da0;
mem_array[4748] = 16'hbdd4;
mem_array[4751] = 16'h547d;
mem_array[4750] = 16'hbf12;
mem_array[4753] = 16'hd84a;
mem_array[4752] = 16'h3f49;
mem_array[4755] = 16'h1582;
mem_array[4754] = 16'h3eef;
mem_array[4757] = 16'h11e3;
mem_array[4756] = 16'h3f52;
mem_array[4759] = 16'h696e;
mem_array[4758] = 16'hbc5b;
mem_array[4761] = 16'hbaf0;
mem_array[4760] = 16'hbca5;
mem_array[4763] = 16'h66c4;
mem_array[4762] = 16'h3d30;
mem_array[4765] = 16'h7c76;
mem_array[4764] = 16'h3e0a;
mem_array[4767] = 16'h5740;
mem_array[4766] = 16'h3eb8;
mem_array[4769] = 16'h7020;
mem_array[4768] = 16'h3f79;
mem_array[4771] = 16'h2776;
mem_array[4770] = 16'hbf92;
mem_array[4773] = 16'hb644;
mem_array[4772] = 16'h3e7e;
mem_array[4775] = 16'h8421;
mem_array[4774] = 16'hbd9c;
mem_array[4777] = 16'h00da;
mem_array[4776] = 16'hbe63;
mem_array[4779] = 16'h8b79;
mem_array[4778] = 16'hbed1;
mem_array[4781] = 16'ha58b;
mem_array[4780] = 16'hbe3a;
mem_array[4783] = 16'h61b6;
mem_array[4782] = 16'h3dc1;
mem_array[4785] = 16'h3525;
mem_array[4784] = 16'hbd4a;
mem_array[4787] = 16'h5515;
mem_array[4786] = 16'h3e17;
mem_array[4789] = 16'h0d69;
mem_array[4788] = 16'h3edc;
mem_array[4791] = 16'h76b5;
mem_array[4790] = 16'h3d45;
mem_array[4793] = 16'hcb84;
mem_array[4792] = 16'hbe7c;
mem_array[4795] = 16'h8590;
mem_array[4794] = 16'hbd9c;
mem_array[4797] = 16'hb3b6;
mem_array[4796] = 16'h3f84;
mem_array[4799] = 16'hc699;
mem_array[4798] = 16'hbe3c;
mem_array[4801] = 16'h0a17;
mem_array[4800] = 16'h3c12;
mem_array[4803] = 16'hb245;
mem_array[4802] = 16'hbd7b;
mem_array[4805] = 16'hb392;
mem_array[4804] = 16'hba3b;
mem_array[4807] = 16'h09e5;
mem_array[4806] = 16'hbdaa;
mem_array[4809] = 16'h6f89;
mem_array[4808] = 16'hbbe3;
mem_array[4811] = 16'h3d15;
mem_array[4810] = 16'hbe50;
mem_array[4813] = 16'h2613;
mem_array[4812] = 16'h3f57;
mem_array[4815] = 16'h8235;
mem_array[4814] = 16'hbb9c;
mem_array[4817] = 16'he0ce;
mem_array[4816] = 16'h3f44;
mem_array[4819] = 16'h3e6b;
mem_array[4818] = 16'hbd14;
mem_array[4821] = 16'h33de;
mem_array[4820] = 16'h3c88;
mem_array[4823] = 16'h02bc;
mem_array[4822] = 16'hbd10;
mem_array[4825] = 16'h314f;
mem_array[4824] = 16'h3dcf;
mem_array[4827] = 16'h40ce;
mem_array[4826] = 16'h3ecc;
mem_array[4829] = 16'h3036;
mem_array[4828] = 16'h3c93;
mem_array[4831] = 16'h08bc;
mem_array[4830] = 16'hbe85;
mem_array[4833] = 16'h23db;
mem_array[4832] = 16'hbd75;
mem_array[4835] = 16'h68f7;
mem_array[4834] = 16'h3d4c;
mem_array[4837] = 16'h85bb;
mem_array[4836] = 16'hbd5f;
mem_array[4839] = 16'h5e10;
mem_array[4838] = 16'hbc78;
mem_array[4841] = 16'he83c;
mem_array[4840] = 16'hbca2;
mem_array[4843] = 16'hbf7e;
mem_array[4842] = 16'hbe9f;
mem_array[4845] = 16'he760;
mem_array[4844] = 16'hbd98;
mem_array[4847] = 16'h3ffe;
mem_array[4846] = 16'hbe9f;
mem_array[4849] = 16'h3e91;
mem_array[4848] = 16'h3e83;
mem_array[4851] = 16'h1a1f;
mem_array[4850] = 16'h3bf3;
mem_array[4853] = 16'h6931;
mem_array[4852] = 16'h3f10;
mem_array[4855] = 16'hebd1;
mem_array[4854] = 16'hbd25;
mem_array[4857] = 16'h28da;
mem_array[4856] = 16'h3f1a;
mem_array[4859] = 16'h88c9;
mem_array[4858] = 16'hbc88;
mem_array[4861] = 16'h758c;
mem_array[4860] = 16'h3daa;
mem_array[4863] = 16'h5dcb;
mem_array[4862] = 16'hbcc0;
mem_array[4865] = 16'h7826;
mem_array[4864] = 16'hbcec;
mem_array[4867] = 16'h3f0a;
mem_array[4866] = 16'h3b70;
mem_array[4869] = 16'h9f57;
mem_array[4868] = 16'hba82;
mem_array[4871] = 16'haa3b;
mem_array[4870] = 16'hbe8d;
mem_array[4873] = 16'hc4bf;
mem_array[4872] = 16'h3f5e;
mem_array[4875] = 16'hdac8;
mem_array[4874] = 16'h3d29;
mem_array[4877] = 16'h4363;
mem_array[4876] = 16'h3f44;
mem_array[4879] = 16'h9f65;
mem_array[4878] = 16'h3c8b;
mem_array[4881] = 16'h698f;
mem_array[4880] = 16'hbdc2;
mem_array[4883] = 16'hda3e;
mem_array[4882] = 16'hbdb0;
mem_array[4885] = 16'h591d;
mem_array[4884] = 16'hbe99;
mem_array[4887] = 16'h5775;
mem_array[4886] = 16'h3f43;
mem_array[4889] = 16'h8f43;
mem_array[4888] = 16'h3df3;
mem_array[4891] = 16'h37ae;
mem_array[4890] = 16'h3d85;
mem_array[4893] = 16'hbf80;
mem_array[4892] = 16'h3ddd;
mem_array[4895] = 16'h80a5;
mem_array[4894] = 16'h3c31;
mem_array[4897] = 16'hac75;
mem_array[4896] = 16'hbdbc;
mem_array[4899] = 16'h7dbe;
mem_array[4898] = 16'hbc96;
mem_array[4901] = 16'ha608;
mem_array[4900] = 16'hbad7;
mem_array[4903] = 16'heb17;
mem_array[4902] = 16'hbe2f;
mem_array[4905] = 16'h416c;
mem_array[4904] = 16'hbe5a;
mem_array[4907] = 16'h4a4a;
mem_array[4906] = 16'hbf5e;
mem_array[4909] = 16'h1176;
mem_array[4908] = 16'h3e3d;
mem_array[4911] = 16'h82ed;
mem_array[4910] = 16'hbda2;
mem_array[4913] = 16'h25f7;
mem_array[4912] = 16'h3f46;
mem_array[4915] = 16'hd70f;
mem_array[4914] = 16'hbda1;
mem_array[4917] = 16'h9ab0;
mem_array[4916] = 16'h3f1f;
mem_array[4919] = 16'h3379;
mem_array[4918] = 16'hbe89;
mem_array[4921] = 16'hfbaf;
mem_array[4920] = 16'hbdb4;
mem_array[4923] = 16'h8a6a;
mem_array[4922] = 16'h3cdc;
mem_array[4925] = 16'h4527;
mem_array[4924] = 16'h3d84;
mem_array[4927] = 16'he838;
mem_array[4926] = 16'h3d98;
mem_array[4929] = 16'h089c;
mem_array[4928] = 16'hbdb8;
mem_array[4931] = 16'h418a;
mem_array[4930] = 16'hbce3;
mem_array[4933] = 16'h07b4;
mem_array[4932] = 16'h3d76;
mem_array[4935] = 16'h8afc;
mem_array[4934] = 16'h3ddd;
mem_array[4937] = 16'h08e9;
mem_array[4936] = 16'hbc9a;
mem_array[4939] = 16'haaf7;
mem_array[4938] = 16'hbde0;
mem_array[4941] = 16'h9b64;
mem_array[4940] = 16'h3dba;
mem_array[4943] = 16'h92d4;
mem_array[4942] = 16'hbca8;
mem_array[4945] = 16'h6482;
mem_array[4944] = 16'hbc08;
mem_array[4947] = 16'h1a0a;
mem_array[4946] = 16'h3cd5;
mem_array[4949] = 16'h8510;
mem_array[4948] = 16'hbcdc;
mem_array[4951] = 16'h5cb3;
mem_array[4950] = 16'h3d21;
mem_array[4953] = 16'h9cde;
mem_array[4952] = 16'h3d8c;
mem_array[4955] = 16'hf247;
mem_array[4954] = 16'h3d4c;
mem_array[4957] = 16'hdd5f;
mem_array[4956] = 16'h3be3;
mem_array[4959] = 16'h3550;
mem_array[4958] = 16'hbdc1;
mem_array[4961] = 16'hfd83;
mem_array[4960] = 16'hbd00;
mem_array[4963] = 16'h4f57;
mem_array[4962] = 16'hbd5c;
mem_array[4965] = 16'hf167;
mem_array[4964] = 16'h3c12;
mem_array[4967] = 16'h4da5;
mem_array[4966] = 16'h3cca;
mem_array[4969] = 16'ha792;
mem_array[4968] = 16'hbcbf;
mem_array[4971] = 16'hdf14;
mem_array[4970] = 16'h3b13;
mem_array[4973] = 16'h885e;
mem_array[4972] = 16'hbbe0;
mem_array[4975] = 16'hd65e;
mem_array[4974] = 16'h3dd5;
mem_array[4977] = 16'h83b3;
mem_array[4976] = 16'h3cac;
mem_array[4979] = 16'h28fc;
mem_array[4978] = 16'hbbb9;
mem_array[4981] = 16'h5b7e;
mem_array[4980] = 16'h3cce;
mem_array[4983] = 16'h5c0f;
mem_array[4982] = 16'h3d10;
mem_array[4985] = 16'h6dbc;
mem_array[4984] = 16'hbbbc;
mem_array[4987] = 16'h8d5c;
mem_array[4986] = 16'h3d4f;
mem_array[4989] = 16'he88e;
mem_array[4988] = 16'hbbc1;
mem_array[4991] = 16'ha0a4;
mem_array[4990] = 16'hbd2a;
mem_array[4993] = 16'hfe54;
mem_array[4992] = 16'h3c6d;
mem_array[4995] = 16'he19a;
mem_array[4994] = 16'hbcf7;
mem_array[4997] = 16'hee8f;
mem_array[4996] = 16'hbd47;
mem_array[4999] = 16'h2383;
mem_array[4998] = 16'hbd3d;
mem_array[5001] = 16'he022;
mem_array[5000] = 16'hbd3c;
mem_array[5003] = 16'h3a69;
mem_array[5002] = 16'h3d7c;
mem_array[5005] = 16'hc200;
mem_array[5004] = 16'h3dac;
mem_array[5007] = 16'h6567;
mem_array[5006] = 16'h3c47;
mem_array[5009] = 16'hca11;
mem_array[5008] = 16'h3cf1;
mem_array[5011] = 16'h2278;
mem_array[5010] = 16'hbd3c;
mem_array[5013] = 16'h2c3b;
mem_array[5012] = 16'h3daf;
mem_array[5015] = 16'hafeb;
mem_array[5014] = 16'hbda9;
mem_array[5017] = 16'hf74f;
mem_array[5016] = 16'h3c73;
mem_array[5019] = 16'h26b3;
mem_array[5018] = 16'h3b9e;
mem_array[5021] = 16'h3dd1;
mem_array[5020] = 16'h3db7;
mem_array[5023] = 16'h4a0d;
mem_array[5022] = 16'h3d52;
mem_array[5025] = 16'hed36;
mem_array[5024] = 16'h3c16;
mem_array[5027] = 16'h364f;
mem_array[5026] = 16'h3d64;
mem_array[5029] = 16'h66eb;
mem_array[5028] = 16'h3dcd;
mem_array[5031] = 16'hd93a;
mem_array[5030] = 16'h3dab;
mem_array[5033] = 16'h6728;
mem_array[5032] = 16'hbc40;
mem_array[5035] = 16'ha8ab;
mem_array[5034] = 16'h3d84;
mem_array[5037] = 16'h0f75;
mem_array[5036] = 16'hbdcf;
mem_array[5039] = 16'h0e81;
mem_array[5038] = 16'h3d69;
mem_array[5041] = 16'h6f6f;
mem_array[5040] = 16'hbdcb;
mem_array[5043] = 16'hdf7e;
mem_array[5042] = 16'h3d44;
mem_array[5045] = 16'h5e50;
mem_array[5044] = 16'h3d41;
mem_array[5047] = 16'h6de1;
mem_array[5046] = 16'hbd4e;
mem_array[5049] = 16'hec2d;
mem_array[5048] = 16'h3ce5;
mem_array[5051] = 16'h181c;
mem_array[5050] = 16'h3969;
mem_array[5053] = 16'hc03a;
mem_array[5052] = 16'hbc07;
mem_array[5055] = 16'h0cf5;
mem_array[5054] = 16'h3cd6;
mem_array[5057] = 16'h80e2;
mem_array[5056] = 16'h3db3;
mem_array[5059] = 16'h7fff;
mem_array[5058] = 16'hbc6e;
mem_array[5061] = 16'h7320;
mem_array[5060] = 16'h3d18;
mem_array[5063] = 16'h03bb;
mem_array[5062] = 16'h3c7d;
mem_array[5065] = 16'hf677;
mem_array[5064] = 16'h3d06;
mem_array[5067] = 16'hecf3;
mem_array[5066] = 16'h3d0f;
mem_array[5069] = 16'h8bca;
mem_array[5068] = 16'hbdd4;
mem_array[5071] = 16'hb170;
mem_array[5070] = 16'hbd80;
mem_array[5073] = 16'hfeff;
mem_array[5072] = 16'h3da9;
mem_array[5075] = 16'h6a9b;
mem_array[5074] = 16'h3d4f;
mem_array[5077] = 16'hf062;
mem_array[5076] = 16'hbcd9;
mem_array[5079] = 16'hbc16;
mem_array[5078] = 16'hbc21;
mem_array[5081] = 16'h8e68;
mem_array[5080] = 16'h3d34;
mem_array[5083] = 16'h39c4;
mem_array[5082] = 16'h3cc7;
mem_array[5085] = 16'h82f0;
mem_array[5084] = 16'h3b41;
mem_array[5087] = 16'h3c09;
mem_array[5086] = 16'h3c20;
mem_array[5089] = 16'h58c8;
mem_array[5088] = 16'h3c8e;
mem_array[5091] = 16'hbd24;
mem_array[5090] = 16'hbd0a;
mem_array[5093] = 16'hc81d;
mem_array[5092] = 16'h3bef;
mem_array[5095] = 16'h5c85;
mem_array[5094] = 16'h3d8d;
mem_array[5097] = 16'h499b;
mem_array[5096] = 16'h3d32;
mem_array[5099] = 16'hac14;
mem_array[5098] = 16'h3d22;
mem_array[5101] = 16'h394f;
mem_array[5100] = 16'h3c56;
mem_array[5103] = 16'h5a31;
mem_array[5102] = 16'h3d80;
mem_array[5105] = 16'he6ec;
mem_array[5104] = 16'h3d4a;
mem_array[5107] = 16'h8007;
mem_array[5106] = 16'h3dda;
mem_array[5109] = 16'hb8d6;
mem_array[5108] = 16'h3d87;
mem_array[5111] = 16'hbb74;
mem_array[5110] = 16'hbc9c;
mem_array[5113] = 16'h253d;
mem_array[5112] = 16'h3caa;
mem_array[5115] = 16'h0e86;
mem_array[5114] = 16'hbd1e;
mem_array[5117] = 16'h2fb7;
mem_array[5116] = 16'hbd0c;
mem_array[5119] = 16'hc46a;
mem_array[5118] = 16'h3d8b;
mem_array[5121] = 16'hfe97;
mem_array[5120] = 16'h3d28;
mem_array[5123] = 16'h8be4;
mem_array[5122] = 16'h3d98;
mem_array[5125] = 16'he586;
mem_array[5124] = 16'h3d45;
mem_array[5127] = 16'h2e66;
mem_array[5126] = 16'h3d61;
mem_array[5129] = 16'h861d;
mem_array[5128] = 16'hbc9f;
mem_array[5131] = 16'h24cb;
mem_array[5130] = 16'h3cf6;
mem_array[5133] = 16'h94cc;
mem_array[5132] = 16'h3d90;
mem_array[5135] = 16'h41ef;
mem_array[5134] = 16'hbd8b;
mem_array[5137] = 16'h4994;
mem_array[5136] = 16'h3a81;
mem_array[5139] = 16'h8c07;
mem_array[5138] = 16'hbccd;
mem_array[5141] = 16'h8c56;
mem_array[5140] = 16'h3d1d;
mem_array[5143] = 16'h29d5;
mem_array[5142] = 16'h3c15;
mem_array[5145] = 16'ha168;
mem_array[5144] = 16'h3d5f;
mem_array[5147] = 16'ha280;
mem_array[5146] = 16'h3d61;
mem_array[5149] = 16'h3483;
mem_array[5148] = 16'hbd7f;
mem_array[5151] = 16'hc3a9;
mem_array[5150] = 16'hbc13;
mem_array[5153] = 16'h62e9;
mem_array[5152] = 16'h3d8d;
mem_array[5155] = 16'h5b8b;
mem_array[5154] = 16'hbcb1;
mem_array[5157] = 16'ha5c6;
mem_array[5156] = 16'hbd94;
mem_array[5159] = 16'h1129;
mem_array[5158] = 16'h3d33;
mem_array[5161] = 16'hbced;
mem_array[5160] = 16'h3ee8;
mem_array[5163] = 16'ha98b;
mem_array[5162] = 16'h3a9f;
mem_array[5165] = 16'h8efa;
mem_array[5164] = 16'h3db9;
mem_array[5167] = 16'h8394;
mem_array[5166] = 16'h3c59;
mem_array[5169] = 16'hafe2;
mem_array[5168] = 16'h3b8c;
mem_array[5171] = 16'h5ff8;
mem_array[5170] = 16'h3d95;
mem_array[5173] = 16'ha75a;
mem_array[5172] = 16'hbd1b;
mem_array[5175] = 16'h2145;
mem_array[5174] = 16'hbe2b;
mem_array[5177] = 16'hca6f;
mem_array[5176] = 16'h3d65;
mem_array[5179] = 16'h67a6;
mem_array[5178] = 16'h3f54;
mem_array[5181] = 16'hd9ad;
mem_array[5180] = 16'h3d8f;
mem_array[5183] = 16'hb8d0;
mem_array[5182] = 16'hbc39;
mem_array[5185] = 16'h08ab;
mem_array[5184] = 16'h3d12;
mem_array[5187] = 16'h6bdf;
mem_array[5186] = 16'h3e05;
mem_array[5189] = 16'h77c2;
mem_array[5188] = 16'h3d8f;
mem_array[5191] = 16'h4827;
mem_array[5190] = 16'h3f21;
mem_array[5193] = 16'ha1bc;
mem_array[5192] = 16'h3d88;
mem_array[5195] = 16'hd378;
mem_array[5194] = 16'hbcb7;
mem_array[5197] = 16'h2a3c;
mem_array[5196] = 16'h3dbd;
mem_array[5199] = 16'hd1c1;
mem_array[5198] = 16'h3bb6;
mem_array[5201] = 16'h0cea;
mem_array[5200] = 16'hbe2f;
mem_array[5203] = 16'h3fce;
mem_array[5202] = 16'hbef7;
mem_array[5205] = 16'h8225;
mem_array[5204] = 16'hbf32;
mem_array[5207] = 16'h03d5;
mem_array[5206] = 16'hbf56;
mem_array[5209] = 16'ha2be;
mem_array[5208] = 16'hbe3c;
mem_array[5211] = 16'h28c5;
mem_array[5210] = 16'h3c9b;
mem_array[5213] = 16'h3e77;
mem_array[5212] = 16'h3e11;
mem_array[5215] = 16'h4e8e;
mem_array[5214] = 16'hbd13;
mem_array[5217] = 16'hdd4f;
mem_array[5216] = 16'h3d0c;
mem_array[5219] = 16'h9ce0;
mem_array[5218] = 16'hbe9e;
mem_array[5221] = 16'h4059;
mem_array[5220] = 16'h3f07;
mem_array[5223] = 16'h2ff4;
mem_array[5222] = 16'hbdc6;
mem_array[5225] = 16'haaa7;
mem_array[5224] = 16'h3cb6;
mem_array[5227] = 16'hb7e6;
mem_array[5226] = 16'h3dd6;
mem_array[5229] = 16'h4712;
mem_array[5228] = 16'h3d9c;
mem_array[5231] = 16'h5509;
mem_array[5230] = 16'h3cff;
mem_array[5233] = 16'he00e;
mem_array[5232] = 16'hbded;
mem_array[5235] = 16'h6ecc;
mem_array[5234] = 16'h3f13;
mem_array[5237] = 16'h647e;
mem_array[5236] = 16'h3da7;
mem_array[5239] = 16'hc5aa;
mem_array[5238] = 16'h3f33;
mem_array[5241] = 16'he923;
mem_array[5240] = 16'hbd6c;
mem_array[5243] = 16'hf725;
mem_array[5242] = 16'hbcf3;
mem_array[5245] = 16'h220b;
mem_array[5244] = 16'h3ea1;
mem_array[5247] = 16'hdd8d;
mem_array[5246] = 16'h3e8e;
mem_array[5249] = 16'hfee0;
mem_array[5248] = 16'hbd17;
mem_array[5251] = 16'h06ac;
mem_array[5250] = 16'hbd63;
mem_array[5253] = 16'h2c25;
mem_array[5252] = 16'hbd88;
mem_array[5255] = 16'h616f;
mem_array[5254] = 16'hbecc;
mem_array[5257] = 16'h08dd;
mem_array[5256] = 16'hbe55;
mem_array[5259] = 16'h15f8;
mem_array[5258] = 16'hbf2c;
mem_array[5261] = 16'hdca0;
mem_array[5260] = 16'hbe52;
mem_array[5263] = 16'h7996;
mem_array[5262] = 16'h3d11;
mem_array[5265] = 16'h9788;
mem_array[5264] = 16'hbf41;
mem_array[5267] = 16'h29cd;
mem_array[5266] = 16'hbebb;
mem_array[5269] = 16'h9454;
mem_array[5268] = 16'hbc2e;
mem_array[5271] = 16'he6a3;
mem_array[5270] = 16'h3d25;
mem_array[5273] = 16'h3deb;
mem_array[5272] = 16'h3f24;
mem_array[5275] = 16'h688f;
mem_array[5274] = 16'h3cb7;
mem_array[5277] = 16'h5768;
mem_array[5276] = 16'h3d57;
mem_array[5279] = 16'ha587;
mem_array[5278] = 16'hbf76;
mem_array[5281] = 16'h1b15;
mem_array[5280] = 16'hbd6b;
mem_array[5283] = 16'h6339;
mem_array[5282] = 16'hbe20;
mem_array[5285] = 16'h561e;
mem_array[5284] = 16'h3e4e;
mem_array[5287] = 16'h0633;
mem_array[5286] = 16'h3ec6;
mem_array[5289] = 16'h1790;
mem_array[5288] = 16'h3d5e;
mem_array[5291] = 16'h8d4e;
mem_array[5290] = 16'h3e09;
mem_array[5293] = 16'h168e;
mem_array[5292] = 16'hbd85;
mem_array[5295] = 16'ha0d7;
mem_array[5294] = 16'h3e85;
mem_array[5297] = 16'h7787;
mem_array[5296] = 16'h3af6;
mem_array[5299] = 16'h306d;
mem_array[5298] = 16'hbd9e;
mem_array[5301] = 16'h93ed;
mem_array[5300] = 16'h3d5e;
mem_array[5303] = 16'he128;
mem_array[5302] = 16'hbd92;
mem_array[5305] = 16'hbe0c;
mem_array[5304] = 16'h3edf;
mem_array[5307] = 16'h00c2;
mem_array[5306] = 16'h3c40;
mem_array[5309] = 16'h5719;
mem_array[5308] = 16'h3e05;
mem_array[5311] = 16'h07d8;
mem_array[5310] = 16'hbf09;
mem_array[5313] = 16'h1df4;
mem_array[5312] = 16'h3e12;
mem_array[5315] = 16'ha073;
mem_array[5314] = 16'hbe24;
mem_array[5317] = 16'h815f;
mem_array[5316] = 16'hbec5;
mem_array[5319] = 16'h9635;
mem_array[5318] = 16'hbf2a;
mem_array[5321] = 16'hafb5;
mem_array[5320] = 16'hbbd1;
mem_array[5323] = 16'h0ba2;
mem_array[5322] = 16'h3e00;
mem_array[5325] = 16'h53f8;
mem_array[5324] = 16'h3d49;
mem_array[5327] = 16'h6df7;
mem_array[5326] = 16'h3f3e;
mem_array[5329] = 16'h3d75;
mem_array[5328] = 16'h3e77;
mem_array[5331] = 16'h4e84;
mem_array[5330] = 16'h3dc8;
mem_array[5333] = 16'h898c;
mem_array[5332] = 16'h3e84;
mem_array[5335] = 16'ha8ed;
mem_array[5334] = 16'hbd29;
mem_array[5337] = 16'hea6f;
mem_array[5336] = 16'h3d70;
mem_array[5339] = 16'hbdaa;
mem_array[5338] = 16'hbe5f;
mem_array[5341] = 16'h0599;
mem_array[5340] = 16'h3cae;
mem_array[5343] = 16'h218b;
mem_array[5342] = 16'hbe27;
mem_array[5345] = 16'hcdc8;
mem_array[5344] = 16'h3dc9;
mem_array[5347] = 16'hd301;
mem_array[5346] = 16'hbeb5;
mem_array[5349] = 16'h1138;
mem_array[5348] = 16'hbea6;
mem_array[5351] = 16'h6cb3;
mem_array[5350] = 16'h3dd6;
mem_array[5353] = 16'h3f97;
mem_array[5352] = 16'h3e6a;
mem_array[5355] = 16'h544e;
mem_array[5354] = 16'hbea0;
mem_array[5357] = 16'h7207;
mem_array[5356] = 16'hbde6;
mem_array[5359] = 16'h00cf;
mem_array[5358] = 16'h3e1a;
mem_array[5361] = 16'hd667;
mem_array[5360] = 16'h3d6c;
mem_array[5363] = 16'h9627;
mem_array[5362] = 16'h3dbf;
mem_array[5365] = 16'hce88;
mem_array[5364] = 16'h3e3d;
mem_array[5367] = 16'h8e13;
mem_array[5366] = 16'h3c7f;
mem_array[5369] = 16'h967b;
mem_array[5368] = 16'h3dae;
mem_array[5371] = 16'hec11;
mem_array[5370] = 16'h3e9f;
mem_array[5373] = 16'he86a;
mem_array[5372] = 16'h3f07;
mem_array[5375] = 16'h9835;
mem_array[5374] = 16'hbee5;
mem_array[5377] = 16'h5ce5;
mem_array[5376] = 16'hbeec;
mem_array[5379] = 16'hf521;
mem_array[5378] = 16'h3e5a;
mem_array[5381] = 16'hb1da;
mem_array[5380] = 16'h3f43;
mem_array[5383] = 16'he484;
mem_array[5382] = 16'h3e6e;
mem_array[5385] = 16'h3003;
mem_array[5384] = 16'hbe33;
mem_array[5387] = 16'hdd41;
mem_array[5386] = 16'h3f12;
mem_array[5389] = 16'hcbb7;
mem_array[5388] = 16'hbee6;
mem_array[5391] = 16'h2334;
mem_array[5390] = 16'h3ddf;
mem_array[5393] = 16'had2e;
mem_array[5392] = 16'h3e61;
mem_array[5395] = 16'h0d18;
mem_array[5394] = 16'h3e49;
mem_array[5397] = 16'hbd61;
mem_array[5396] = 16'h3d99;
mem_array[5399] = 16'h48c1;
mem_array[5398] = 16'hbc00;
mem_array[5401] = 16'h0f07;
mem_array[5400] = 16'h3cdd;
mem_array[5403] = 16'hb0a6;
mem_array[5402] = 16'hbd90;
mem_array[5405] = 16'h9f98;
mem_array[5404] = 16'h3ed4;
mem_array[5407] = 16'hbc1a;
mem_array[5406] = 16'hbf5a;
mem_array[5409] = 16'h39e2;
mem_array[5408] = 16'hbdbc;
mem_array[5411] = 16'h7f31;
mem_array[5410] = 16'h3d8b;
mem_array[5413] = 16'hfd0d;
mem_array[5412] = 16'h3f0d;
mem_array[5415] = 16'hdd64;
mem_array[5414] = 16'h3ec6;
mem_array[5417] = 16'h3517;
mem_array[5416] = 16'h3e4e;
mem_array[5419] = 16'h4cab;
mem_array[5418] = 16'h3ed6;
mem_array[5421] = 16'h8b24;
mem_array[5420] = 16'h3d35;
mem_array[5423] = 16'h5f2b;
mem_array[5422] = 16'hbc32;
mem_array[5425] = 16'hf8f3;
mem_array[5424] = 16'h3f0f;
mem_array[5427] = 16'h23c3;
mem_array[5426] = 16'h3f04;
mem_array[5429] = 16'h8cb3;
mem_array[5428] = 16'h3db4;
mem_array[5431] = 16'hf20b;
mem_array[5430] = 16'hbf39;
mem_array[5433] = 16'h4459;
mem_array[5432] = 16'h3f94;
mem_array[5435] = 16'ha449;
mem_array[5434] = 16'hbf3c;
mem_array[5437] = 16'h4ef5;
mem_array[5436] = 16'hbf25;
mem_array[5439] = 16'h60d6;
mem_array[5438] = 16'h3ed6;
mem_array[5441] = 16'h81f9;
mem_array[5440] = 16'h3e51;
mem_array[5443] = 16'h75b4;
mem_array[5442] = 16'h3ea2;
mem_array[5445] = 16'h710a;
mem_array[5444] = 16'hbe98;
mem_array[5447] = 16'ha4fc;
mem_array[5446] = 16'h3f60;
mem_array[5449] = 16'heff5;
mem_array[5448] = 16'hbb04;
mem_array[5451] = 16'h8c02;
mem_array[5450] = 16'hbc5b;
mem_array[5453] = 16'h2f1a;
mem_array[5452] = 16'hbe5f;
mem_array[5455] = 16'h28f5;
mem_array[5454] = 16'hbc52;
mem_array[5457] = 16'h9527;
mem_array[5456] = 16'h3f0a;
mem_array[5459] = 16'hbec6;
mem_array[5458] = 16'hbf0d;
mem_array[5461] = 16'h7d5e;
mem_array[5460] = 16'h3f40;
mem_array[5463] = 16'h0217;
mem_array[5462] = 16'h3d25;
mem_array[5465] = 16'h2159;
mem_array[5464] = 16'h3f38;
mem_array[5467] = 16'h6582;
mem_array[5466] = 16'hbec2;
mem_array[5469] = 16'hd5e2;
mem_array[5468] = 16'hbd9d;
mem_array[5471] = 16'h682c;
mem_array[5470] = 16'h3e32;
mem_array[5473] = 16'hc3bd;
mem_array[5472] = 16'h3f51;
mem_array[5475] = 16'h3a93;
mem_array[5474] = 16'h3f90;
mem_array[5477] = 16'hf09f;
mem_array[5476] = 16'h3ea6;
mem_array[5479] = 16'hd073;
mem_array[5478] = 16'hbeaa;
mem_array[5481] = 16'h67ba;
mem_array[5480] = 16'h3d99;
mem_array[5483] = 16'h4d0c;
mem_array[5482] = 16'hbca5;
mem_array[5485] = 16'hbf2c;
mem_array[5484] = 16'h3e91;
mem_array[5487] = 16'h066e;
mem_array[5486] = 16'h3fc2;
mem_array[5489] = 16'h3914;
mem_array[5488] = 16'h3ed7;
mem_array[5491] = 16'hf59a;
mem_array[5490] = 16'hbf03;
mem_array[5493] = 16'he812;
mem_array[5492] = 16'h3e1c;
mem_array[5495] = 16'h4427;
mem_array[5494] = 16'hbf82;
mem_array[5497] = 16'hd849;
mem_array[5496] = 16'hbf69;
mem_array[5499] = 16'h8a5d;
mem_array[5498] = 16'hbeb6;
mem_array[5501] = 16'hb2a3;
mem_array[5500] = 16'h3e58;
mem_array[5503] = 16'he808;
mem_array[5502] = 16'h3eb5;
mem_array[5505] = 16'hfa20;
mem_array[5504] = 16'hbf1e;
mem_array[5507] = 16'hd5c6;
mem_array[5506] = 16'h3f03;
mem_array[5509] = 16'h149c;
mem_array[5508] = 16'h3f02;
mem_array[5511] = 16'hf909;
mem_array[5510] = 16'h3ea9;
mem_array[5513] = 16'h416c;
mem_array[5512] = 16'h3ee0;
mem_array[5515] = 16'h12ea;
mem_array[5514] = 16'h3ea1;
mem_array[5517] = 16'h8d49;
mem_array[5516] = 16'h3e83;
mem_array[5519] = 16'ha517;
mem_array[5518] = 16'hbf3b;
mem_array[5521] = 16'hbb0f;
mem_array[5520] = 16'h3f1a;
mem_array[5523] = 16'hcebc;
mem_array[5522] = 16'hbdb5;
mem_array[5525] = 16'h89a0;
mem_array[5524] = 16'hbe49;
mem_array[5527] = 16'h5b8d;
mem_array[5526] = 16'hbf85;
mem_array[5529] = 16'ha8df;
mem_array[5528] = 16'h3f37;
mem_array[5531] = 16'h5b09;
mem_array[5530] = 16'hbf1a;
mem_array[5533] = 16'hc827;
mem_array[5532] = 16'h3ef1;
mem_array[5535] = 16'h6012;
mem_array[5534] = 16'h3f1a;
mem_array[5537] = 16'hfc51;
mem_array[5536] = 16'hbe31;
mem_array[5539] = 16'hfcf4;
mem_array[5538] = 16'hbe84;
mem_array[5541] = 16'hd007;
mem_array[5540] = 16'hbdad;
mem_array[5543] = 16'hde5d;
mem_array[5542] = 16'hbd25;
mem_array[5545] = 16'h8997;
mem_array[5544] = 16'h3d39;
mem_array[5547] = 16'h86fc;
mem_array[5546] = 16'h3ea1;
mem_array[5549] = 16'ha7b1;
mem_array[5548] = 16'h3df1;
mem_array[5551] = 16'h634c;
mem_array[5550] = 16'hbdb2;
mem_array[5553] = 16'h399d;
mem_array[5552] = 16'hbd2d;
mem_array[5555] = 16'h63bc;
mem_array[5554] = 16'hbf47;
mem_array[5557] = 16'h3afb;
mem_array[5556] = 16'hbfa3;
mem_array[5559] = 16'hd1bb;
mem_array[5558] = 16'hbeba;
mem_array[5561] = 16'h716f;
mem_array[5560] = 16'hbf1d;
mem_array[5563] = 16'h1814;
mem_array[5562] = 16'h3f7d;
mem_array[5565] = 16'h19cd;
mem_array[5564] = 16'h3e8f;
mem_array[5567] = 16'hd037;
mem_array[5566] = 16'h3f9d;
mem_array[5569] = 16'he22a;
mem_array[5568] = 16'h3dae;
mem_array[5571] = 16'h9d89;
mem_array[5570] = 16'h3d80;
mem_array[5573] = 16'h948d;
mem_array[5572] = 16'h3f42;
mem_array[5575] = 16'habc1;
mem_array[5574] = 16'h3f25;
mem_array[5577] = 16'hea6a;
mem_array[5576] = 16'h3d96;
mem_array[5579] = 16'h5260;
mem_array[5578] = 16'hbe9b;
mem_array[5581] = 16'h77c1;
mem_array[5580] = 16'h3f27;
mem_array[5583] = 16'h8220;
mem_array[5582] = 16'hbec5;
mem_array[5585] = 16'h748e;
mem_array[5584] = 16'h3f05;
mem_array[5587] = 16'h882a;
mem_array[5586] = 16'hbf57;
mem_array[5589] = 16'h6635;
mem_array[5588] = 16'h3f47;
mem_array[5591] = 16'h8882;
mem_array[5590] = 16'hbfdb;
mem_array[5593] = 16'hbb09;
mem_array[5592] = 16'h3e94;
mem_array[5595] = 16'h458d;
mem_array[5594] = 16'h3f4c;
mem_array[5597] = 16'ha403;
mem_array[5596] = 16'h3dc8;
mem_array[5599] = 16'h1076;
mem_array[5598] = 16'h3f0d;
mem_array[5601] = 16'h4f75;
mem_array[5600] = 16'hbd42;
mem_array[5603] = 16'h2d41;
mem_array[5602] = 16'h3dac;
mem_array[5605] = 16'h63ef;
mem_array[5604] = 16'h3ec7;
mem_array[5607] = 16'hc983;
mem_array[5606] = 16'h3f3b;
mem_array[5609] = 16'h8f69;
mem_array[5608] = 16'h3f05;
mem_array[5611] = 16'h333a;
mem_array[5610] = 16'h3ea4;
mem_array[5613] = 16'hc538;
mem_array[5612] = 16'h3f15;
mem_array[5615] = 16'h01ee;
mem_array[5614] = 16'hbf03;
mem_array[5617] = 16'he26d;
mem_array[5616] = 16'hbfb1;
mem_array[5619] = 16'hdb79;
mem_array[5618] = 16'hbe8e;
mem_array[5621] = 16'h2f49;
mem_array[5620] = 16'hbeee;
mem_array[5623] = 16'h537f;
mem_array[5622] = 16'h3f4c;
mem_array[5625] = 16'h16ef;
mem_array[5624] = 16'hbf25;
mem_array[5627] = 16'h537b;
mem_array[5626] = 16'h3fbf;
mem_array[5629] = 16'h89e4;
mem_array[5628] = 16'h3cbc;
mem_array[5631] = 16'ha825;
mem_array[5630] = 16'hbd8c;
mem_array[5633] = 16'h68a7;
mem_array[5632] = 16'h3eb1;
mem_array[5635] = 16'h6ed1;
mem_array[5634] = 16'hbe06;
mem_array[5637] = 16'hd9f9;
mem_array[5636] = 16'h3f5f;
mem_array[5639] = 16'h9b4a;
mem_array[5638] = 16'hbd98;
mem_array[5641] = 16'h9037;
mem_array[5640] = 16'h3f34;
mem_array[5643] = 16'hf223;
mem_array[5642] = 16'hbf09;
mem_array[5645] = 16'hc96f;
mem_array[5644] = 16'h3f09;
mem_array[5647] = 16'hccd3;
mem_array[5646] = 16'hbe90;
mem_array[5649] = 16'hfcc5;
mem_array[5648] = 16'hbe9e;
mem_array[5651] = 16'he8b7;
mem_array[5650] = 16'hbfb7;
mem_array[5653] = 16'hb151;
mem_array[5652] = 16'h3f3e;
mem_array[5655] = 16'h88a6;
mem_array[5654] = 16'h3f1f;
mem_array[5657] = 16'h80dc;
mem_array[5656] = 16'hbec7;
mem_array[5659] = 16'hfbcf;
mem_array[5658] = 16'h3ed2;
mem_array[5661] = 16'h1a73;
mem_array[5660] = 16'h3da4;
mem_array[5663] = 16'h2d6b;
mem_array[5662] = 16'hbd32;
mem_array[5665] = 16'hc813;
mem_array[5664] = 16'h3e51;
mem_array[5667] = 16'h00e6;
mem_array[5666] = 16'h3ea7;
mem_array[5669] = 16'h36e3;
mem_array[5668] = 16'h3f18;
mem_array[5671] = 16'h0734;
mem_array[5670] = 16'h3e84;
mem_array[5673] = 16'h769b;
mem_array[5672] = 16'h3e36;
mem_array[5675] = 16'h7e28;
mem_array[5674] = 16'hbeab;
mem_array[5677] = 16'h40f1;
mem_array[5676] = 16'hbfea;
mem_array[5679] = 16'hb397;
mem_array[5678] = 16'h3e70;
mem_array[5681] = 16'h5978;
mem_array[5680] = 16'hbf14;
mem_array[5683] = 16'h4d73;
mem_array[5682] = 16'h3f22;
mem_array[5685] = 16'he4ad;
mem_array[5684] = 16'hbf75;
mem_array[5687] = 16'h21fd;
mem_array[5686] = 16'h3fa2;
mem_array[5689] = 16'h9640;
mem_array[5688] = 16'hbf23;
mem_array[5691] = 16'h9b1f;
mem_array[5690] = 16'hbf05;
mem_array[5693] = 16'h2c6b;
mem_array[5692] = 16'h3e64;
mem_array[5695] = 16'h2f7a;
mem_array[5694] = 16'hbef5;
mem_array[5697] = 16'h81be;
mem_array[5696] = 16'h3f98;
mem_array[5699] = 16'h51d2;
mem_array[5698] = 16'h3e90;
mem_array[5701] = 16'h293d;
mem_array[5700] = 16'h3e2c;
mem_array[5703] = 16'h81b6;
mem_array[5702] = 16'hbf3f;
mem_array[5705] = 16'h2684;
mem_array[5704] = 16'h3db8;
mem_array[5707] = 16'h01ff;
mem_array[5706] = 16'hbe05;
mem_array[5709] = 16'hbb82;
mem_array[5708] = 16'h3ba0;
mem_array[5711] = 16'h43c0;
mem_array[5710] = 16'hbfad;
mem_array[5713] = 16'h7ea5;
mem_array[5712] = 16'h3f1c;
mem_array[5715] = 16'h5619;
mem_array[5714] = 16'h3f23;
mem_array[5717] = 16'hae10;
mem_array[5716] = 16'hbe0f;
mem_array[5719] = 16'haa3b;
mem_array[5718] = 16'hbeab;
mem_array[5721] = 16'hdc48;
mem_array[5720] = 16'h3be3;
mem_array[5723] = 16'h7b64;
mem_array[5722] = 16'h3cc0;
mem_array[5725] = 16'h1d43;
mem_array[5724] = 16'h3ea2;
mem_array[5727] = 16'hcc82;
mem_array[5726] = 16'h3eb0;
mem_array[5729] = 16'h57f4;
mem_array[5728] = 16'h3f99;
mem_array[5731] = 16'hb510;
mem_array[5730] = 16'h3f41;
mem_array[5733] = 16'h722f;
mem_array[5732] = 16'h3e44;
mem_array[5735] = 16'h39b1;
mem_array[5734] = 16'hbe60;
mem_array[5737] = 16'h1fd9;
mem_array[5736] = 16'hbff8;
mem_array[5739] = 16'h1b42;
mem_array[5738] = 16'h3e1e;
mem_array[5741] = 16'hf526;
mem_array[5740] = 16'h3c94;
mem_array[5743] = 16'h45af;
mem_array[5742] = 16'h3f12;
mem_array[5745] = 16'hf0c9;
mem_array[5744] = 16'hbf1d;
mem_array[5747] = 16'h6efe;
mem_array[5746] = 16'h3f97;
mem_array[5749] = 16'hdaa7;
mem_array[5748] = 16'hbeb6;
mem_array[5751] = 16'hd1c5;
mem_array[5750] = 16'hbeb2;
mem_array[5753] = 16'h3afd;
mem_array[5752] = 16'h3f31;
mem_array[5755] = 16'hc659;
mem_array[5754] = 16'hbd80;
mem_array[5757] = 16'h4128;
mem_array[5756] = 16'h3f51;
mem_array[5759] = 16'h7bdb;
mem_array[5758] = 16'h3ea2;
mem_array[5761] = 16'h906c;
mem_array[5760] = 16'hbe91;
mem_array[5763] = 16'h2b75;
mem_array[5762] = 16'hbe9f;
mem_array[5765] = 16'hed97;
mem_array[5764] = 16'hbf1a;
mem_array[5767] = 16'h3b32;
mem_array[5766] = 16'hbf23;
mem_array[5769] = 16'h964f;
mem_array[5768] = 16'h3eb7;
mem_array[5771] = 16'h5af0;
mem_array[5770] = 16'h3dcc;
mem_array[5773] = 16'hb8db;
mem_array[5772] = 16'h3f86;
mem_array[5775] = 16'h6a1d;
mem_array[5774] = 16'h3f9a;
mem_array[5777] = 16'h5075;
mem_array[5776] = 16'hbf15;
mem_array[5779] = 16'h415c;
mem_array[5778] = 16'h3f62;
mem_array[5781] = 16'h6d6e;
mem_array[5780] = 16'hbdbc;
mem_array[5783] = 16'h3ef1;
mem_array[5782] = 16'h3cca;
mem_array[5785] = 16'h2b29;
mem_array[5784] = 16'hbc5d;
mem_array[5787] = 16'ha610;
mem_array[5786] = 16'hbde1;
mem_array[5789] = 16'ha429;
mem_array[5788] = 16'h3d92;
mem_array[5791] = 16'h8e24;
mem_array[5790] = 16'h3ee5;
mem_array[5793] = 16'h9827;
mem_array[5792] = 16'h3f22;
mem_array[5795] = 16'h250f;
mem_array[5794] = 16'hbd71;
mem_array[5797] = 16'h81f3;
mem_array[5796] = 16'hbf95;
mem_array[5799] = 16'h6a05;
mem_array[5798] = 16'h3d93;
mem_array[5801] = 16'h6cea;
mem_array[5800] = 16'hbf00;
mem_array[5803] = 16'h86cd;
mem_array[5802] = 16'h3e9c;
mem_array[5805] = 16'hed24;
mem_array[5804] = 16'hbf7c;
mem_array[5807] = 16'hf860;
mem_array[5806] = 16'h3f5e;
mem_array[5809] = 16'hc273;
mem_array[5808] = 16'hbf0f;
mem_array[5811] = 16'h8459;
mem_array[5810] = 16'hbec5;
mem_array[5813] = 16'h844f;
mem_array[5812] = 16'h3f52;
mem_array[5815] = 16'h68f9;
mem_array[5814] = 16'h3e15;
mem_array[5817] = 16'ha4bf;
mem_array[5816] = 16'h3df3;
mem_array[5819] = 16'h4cd8;
mem_array[5818] = 16'hbe8a;
mem_array[5821] = 16'h7d44;
mem_array[5820] = 16'hbf5a;
mem_array[5823] = 16'h6b4b;
mem_array[5822] = 16'hbf02;
mem_array[5825] = 16'h239d;
mem_array[5824] = 16'hbeb1;
mem_array[5827] = 16'hc6b6;
mem_array[5826] = 16'hbf38;
mem_array[5829] = 16'he927;
mem_array[5828] = 16'h3e13;
mem_array[5831] = 16'h8b92;
mem_array[5830] = 16'h3f38;
mem_array[5833] = 16'h1e7f;
mem_array[5832] = 16'h3ebb;
mem_array[5835] = 16'h5d1a;
mem_array[5834] = 16'h3f63;
mem_array[5837] = 16'h959d;
mem_array[5836] = 16'hbf70;
mem_array[5839] = 16'h64fa;
mem_array[5838] = 16'h3f17;
mem_array[5841] = 16'h7aac;
mem_array[5840] = 16'h3c73;
mem_array[5843] = 16'hc306;
mem_array[5842] = 16'h3d22;
mem_array[5845] = 16'hd9a1;
mem_array[5844] = 16'h3f27;
mem_array[5847] = 16'h503e;
mem_array[5846] = 16'h3e82;
mem_array[5849] = 16'he9e5;
mem_array[5848] = 16'h3ed4;
mem_array[5851] = 16'ha5a0;
mem_array[5850] = 16'h3e80;
mem_array[5853] = 16'h4c9a;
mem_array[5852] = 16'h3f0b;
mem_array[5855] = 16'h52cb;
mem_array[5854] = 16'h3dd3;
mem_array[5857] = 16'hf51f;
mem_array[5856] = 16'hc040;
mem_array[5859] = 16'hdbe5;
mem_array[5858] = 16'h3c23;
mem_array[5861] = 16'hffd7;
mem_array[5860] = 16'hbf6f;
mem_array[5863] = 16'h1f53;
mem_array[5862] = 16'h3e16;
mem_array[5865] = 16'hb7b9;
mem_array[5864] = 16'hbee5;
mem_array[5867] = 16'h47e9;
mem_array[5866] = 16'h3f2e;
mem_array[5869] = 16'hbda6;
mem_array[5868] = 16'hbed2;
mem_array[5871] = 16'h11cd;
mem_array[5870] = 16'hbf02;
mem_array[5873] = 16'hda5b;
mem_array[5872] = 16'h3e63;
mem_array[5875] = 16'h80fd;
mem_array[5874] = 16'hbeb1;
mem_array[5877] = 16'he974;
mem_array[5876] = 16'h3ed9;
mem_array[5879] = 16'hfc20;
mem_array[5878] = 16'hbee8;
mem_array[5881] = 16'h716d;
mem_array[5880] = 16'hbff4;
mem_array[5883] = 16'h6d63;
mem_array[5882] = 16'hbf2b;
mem_array[5885] = 16'h1c1a;
mem_array[5884] = 16'hbf05;
mem_array[5887] = 16'haa34;
mem_array[5886] = 16'h3e1e;
mem_array[5889] = 16'hd760;
mem_array[5888] = 16'h3ee4;
mem_array[5891] = 16'hd95e;
mem_array[5890] = 16'h3cfd;
mem_array[5893] = 16'hb70b;
mem_array[5892] = 16'h3e85;
mem_array[5895] = 16'h1fa6;
mem_array[5894] = 16'h3f6c;
mem_array[5897] = 16'hdd41;
mem_array[5896] = 16'hbee7;
mem_array[5899] = 16'h8825;
mem_array[5898] = 16'h3d1d;
mem_array[5901] = 16'h8ce7;
mem_array[5900] = 16'h3c7e;
mem_array[5903] = 16'h9b1d;
mem_array[5902] = 16'hbd14;
mem_array[5905] = 16'hcd87;
mem_array[5904] = 16'h3df9;
mem_array[5907] = 16'he0db;
mem_array[5906] = 16'hbe64;
mem_array[5909] = 16'h00e3;
mem_array[5908] = 16'hbe5b;
mem_array[5911] = 16'hb377;
mem_array[5910] = 16'h3eb5;
mem_array[5913] = 16'h4e04;
mem_array[5912] = 16'h3ee8;
mem_array[5915] = 16'h19e0;
mem_array[5914] = 16'hbe95;
mem_array[5917] = 16'h633a;
mem_array[5916] = 16'hbf73;
mem_array[5919] = 16'h87bf;
mem_array[5918] = 16'hbd8c;
mem_array[5921] = 16'hb809;
mem_array[5920] = 16'h3c9b;
mem_array[5923] = 16'h01d6;
mem_array[5922] = 16'h3e80;
mem_array[5925] = 16'h13d8;
mem_array[5924] = 16'hbd28;
mem_array[5927] = 16'h6cf3;
mem_array[5926] = 16'h3f54;
mem_array[5929] = 16'h80b0;
mem_array[5928] = 16'hbe12;
mem_array[5931] = 16'hfd5f;
mem_array[5930] = 16'h3efe;
mem_array[5933] = 16'hb6d2;
mem_array[5932] = 16'hbd4e;
mem_array[5935] = 16'h97b4;
mem_array[5934] = 16'hbda6;
mem_array[5937] = 16'h8b67;
mem_array[5936] = 16'h3f45;
mem_array[5939] = 16'he6d3;
mem_array[5938] = 16'hbe3f;
mem_array[5941] = 16'h5aa9;
mem_array[5940] = 16'hbf92;
mem_array[5943] = 16'he828;
mem_array[5942] = 16'h3eea;
mem_array[5945] = 16'h2ec6;
mem_array[5944] = 16'hbe34;
mem_array[5947] = 16'h3ad0;
mem_array[5946] = 16'hbe72;
mem_array[5949] = 16'h58ed;
mem_array[5948] = 16'h3ef4;
mem_array[5951] = 16'h986e;
mem_array[5950] = 16'h3eca;
mem_array[5953] = 16'h2bb8;
mem_array[5952] = 16'hbeee;
mem_array[5955] = 16'h2dbb;
mem_array[5954] = 16'h3f43;
mem_array[5957] = 16'h45ea;
mem_array[5956] = 16'hbe9b;
mem_array[5959] = 16'h05c1;
mem_array[5958] = 16'h3f4a;
mem_array[5961] = 16'h7605;
mem_array[5960] = 16'hbd95;
mem_array[5963] = 16'ha816;
mem_array[5962] = 16'hbce8;
mem_array[5965] = 16'h46bb;
mem_array[5964] = 16'h3b78;
mem_array[5967] = 16'h1978;
mem_array[5966] = 16'hbe03;
mem_array[5969] = 16'h2556;
mem_array[5968] = 16'hbeb8;
mem_array[5971] = 16'h6a60;
mem_array[5970] = 16'h3ed7;
mem_array[5973] = 16'h7674;
mem_array[5972] = 16'h3e9f;
mem_array[5975] = 16'h9c41;
mem_array[5974] = 16'hbf26;
mem_array[5977] = 16'h6316;
mem_array[5976] = 16'hbfb5;
mem_array[5979] = 16'hf3f6;
mem_array[5978] = 16'hbd78;
mem_array[5981] = 16'h250c;
mem_array[5980] = 16'hbf93;
mem_array[5983] = 16'h08ed;
mem_array[5982] = 16'h3d92;
mem_array[5985] = 16'hdc28;
mem_array[5984] = 16'hbe41;
mem_array[5987] = 16'h10d0;
mem_array[5986] = 16'h3f33;
mem_array[5989] = 16'h5a44;
mem_array[5988] = 16'hbe1c;
mem_array[5991] = 16'hfd00;
mem_array[5990] = 16'h3eb0;
mem_array[5993] = 16'h777e;
mem_array[5992] = 16'h3dac;
mem_array[5995] = 16'haf8a;
mem_array[5994] = 16'h3e30;
mem_array[5997] = 16'h840b;
mem_array[5996] = 16'h3f13;
mem_array[5999] = 16'h316d;
mem_array[5998] = 16'hbe80;
mem_array[6001] = 16'h0ea5;
mem_array[6000] = 16'hbead;
mem_array[6003] = 16'haabe;
mem_array[6002] = 16'h3e81;
mem_array[6005] = 16'h777d;
mem_array[6004] = 16'hbf25;
mem_array[6007] = 16'h868b;
mem_array[6006] = 16'h3eb6;
mem_array[6009] = 16'hdc0a;
mem_array[6008] = 16'h3efb;
mem_array[6011] = 16'h151a;
mem_array[6010] = 16'h3e0c;
mem_array[6013] = 16'h04bd;
mem_array[6012] = 16'hbf18;
mem_array[6015] = 16'h553c;
mem_array[6014] = 16'h3f51;
mem_array[6017] = 16'h4971;
mem_array[6016] = 16'h3ea4;
mem_array[6019] = 16'h7dc8;
mem_array[6018] = 16'h3f15;
mem_array[6021] = 16'h63ec;
mem_array[6020] = 16'h3d83;
mem_array[6023] = 16'h1870;
mem_array[6022] = 16'h3d72;
mem_array[6025] = 16'he112;
mem_array[6024] = 16'h3e40;
mem_array[6027] = 16'hf4f1;
mem_array[6026] = 16'hbdb0;
mem_array[6029] = 16'h7866;
mem_array[6028] = 16'hbb13;
mem_array[6031] = 16'h3a7a;
mem_array[6030] = 16'h3e77;
mem_array[6033] = 16'hfb75;
mem_array[6032] = 16'h3e24;
mem_array[6035] = 16'h205a;
mem_array[6034] = 16'hbf09;
mem_array[6037] = 16'h8e7a;
mem_array[6036] = 16'hbf28;
mem_array[6039] = 16'h39d9;
mem_array[6038] = 16'h3b49;
mem_array[6041] = 16'haa77;
mem_array[6040] = 16'hbfbc;
mem_array[6043] = 16'h21c7;
mem_array[6042] = 16'h3ea9;
mem_array[6045] = 16'h6de2;
mem_array[6044] = 16'h3ddf;
mem_array[6047] = 16'hdfab;
mem_array[6046] = 16'h3f2a;
mem_array[6049] = 16'h447c;
mem_array[6048] = 16'h3da5;
mem_array[6051] = 16'hf679;
mem_array[6050] = 16'hbe0a;
mem_array[6053] = 16'hc10b;
mem_array[6052] = 16'hbe96;
mem_array[6055] = 16'h437c;
mem_array[6054] = 16'h3f13;
mem_array[6057] = 16'h63fa;
mem_array[6056] = 16'h3f19;
mem_array[6059] = 16'h8223;
mem_array[6058] = 16'hbe2f;
mem_array[6061] = 16'h4009;
mem_array[6060] = 16'h3e06;
mem_array[6063] = 16'heb81;
mem_array[6062] = 16'hbcbe;
mem_array[6065] = 16'hb614;
mem_array[6064] = 16'hbf2e;
mem_array[6067] = 16'he3f1;
mem_array[6066] = 16'hbee1;
mem_array[6069] = 16'he6bf;
mem_array[6068] = 16'h3dc0;
mem_array[6071] = 16'haaef;
mem_array[6070] = 16'h3eba;
mem_array[6073] = 16'hb21b;
mem_array[6072] = 16'h3ed2;
mem_array[6075] = 16'h9a0e;
mem_array[6074] = 16'h3e56;
mem_array[6077] = 16'hffe6;
mem_array[6076] = 16'h3e93;
mem_array[6079] = 16'h8f08;
mem_array[6078] = 16'h3e67;
mem_array[6081] = 16'h5bdc;
mem_array[6080] = 16'hbda4;
mem_array[6083] = 16'hd136;
mem_array[6082] = 16'h3d25;
mem_array[6085] = 16'h6c73;
mem_array[6084] = 16'h3e5d;
mem_array[6087] = 16'h42a5;
mem_array[6086] = 16'h3c6b;
mem_array[6089] = 16'he7b9;
mem_array[6088] = 16'h3e94;
mem_array[6091] = 16'h5c8e;
mem_array[6090] = 16'h3eca;
mem_array[6093] = 16'h8a8c;
mem_array[6092] = 16'h3dca;
mem_array[6095] = 16'h5aef;
mem_array[6094] = 16'hbec4;
mem_array[6097] = 16'h371f;
mem_array[6096] = 16'hbdb5;
mem_array[6099] = 16'hbbc4;
mem_array[6098] = 16'hbd9d;
mem_array[6101] = 16'h6edf;
mem_array[6100] = 16'hbecc;
mem_array[6103] = 16'h1675;
mem_array[6102] = 16'h3dd8;
mem_array[6105] = 16'hc42e;
mem_array[6104] = 16'hbd9d;
mem_array[6107] = 16'h01ba;
mem_array[6106] = 16'h3f25;
mem_array[6109] = 16'h7f73;
mem_array[6108] = 16'h3e8c;
mem_array[6111] = 16'he705;
mem_array[6110] = 16'hbe9f;
mem_array[6113] = 16'h48d2;
mem_array[6112] = 16'hbe15;
mem_array[6115] = 16'hae49;
mem_array[6114] = 16'h3ee0;
mem_array[6117] = 16'h18e1;
mem_array[6116] = 16'h3f72;
mem_array[6119] = 16'he12b;
mem_array[6118] = 16'hbe31;
mem_array[6121] = 16'hc418;
mem_array[6120] = 16'h3eb4;
mem_array[6123] = 16'hf27f;
mem_array[6122] = 16'hbdf4;
mem_array[6125] = 16'hfa9c;
mem_array[6124] = 16'hbf90;
mem_array[6127] = 16'h4516;
mem_array[6126] = 16'hbf24;
mem_array[6129] = 16'h08b6;
mem_array[6128] = 16'h3d89;
mem_array[6131] = 16'h5893;
mem_array[6130] = 16'h3f3d;
mem_array[6133] = 16'h2b2d;
mem_array[6132] = 16'h3bc5;
mem_array[6135] = 16'h481f;
mem_array[6134] = 16'h3efe;
mem_array[6137] = 16'h65fc;
mem_array[6136] = 16'hbe07;
mem_array[6139] = 16'h76c6;
mem_array[6138] = 16'h3e36;
mem_array[6141] = 16'h7a04;
mem_array[6140] = 16'h3db0;
mem_array[6143] = 16'h021c;
mem_array[6142] = 16'hbbee;
mem_array[6145] = 16'hbf9b;
mem_array[6144] = 16'hbdc2;
mem_array[6147] = 16'hf91b;
mem_array[6146] = 16'hbcbf;
mem_array[6149] = 16'h5814;
mem_array[6148] = 16'h3f07;
mem_array[6151] = 16'ha85e;
mem_array[6150] = 16'h3da5;
mem_array[6153] = 16'h376f;
mem_array[6152] = 16'hbd00;
mem_array[6155] = 16'haffb;
mem_array[6154] = 16'hbec6;
mem_array[6157] = 16'h0f92;
mem_array[6156] = 16'hbeee;
mem_array[6159] = 16'hb7da;
mem_array[6158] = 16'hbde6;
mem_array[6161] = 16'hf0fa;
mem_array[6160] = 16'hbf3e;
mem_array[6163] = 16'hde99;
mem_array[6162] = 16'h3e8e;
mem_array[6165] = 16'h1058;
mem_array[6164] = 16'hbe36;
mem_array[6167] = 16'habc9;
mem_array[6166] = 16'h3f50;
mem_array[6169] = 16'h5c5e;
mem_array[6168] = 16'h3ef5;
mem_array[6171] = 16'hed9e;
mem_array[6170] = 16'hbe99;
mem_array[6173] = 16'haca5;
mem_array[6172] = 16'h3d70;
mem_array[6175] = 16'hdd6d;
mem_array[6174] = 16'h3f2c;
mem_array[6177] = 16'h52f6;
mem_array[6176] = 16'h3ede;
mem_array[6179] = 16'h0b99;
mem_array[6178] = 16'hbe60;
mem_array[6181] = 16'hbf5a;
mem_array[6180] = 16'h3e78;
mem_array[6183] = 16'h5f7b;
mem_array[6182] = 16'hbdae;
mem_array[6185] = 16'h1ec7;
mem_array[6184] = 16'hbecf;
mem_array[6187] = 16'hf4fe;
mem_array[6186] = 16'hbf33;
mem_array[6189] = 16'h94ae;
mem_array[6188] = 16'h3ee1;
mem_array[6191] = 16'h9784;
mem_array[6190] = 16'h3dd0;
mem_array[6193] = 16'hdf09;
mem_array[6192] = 16'hbe1c;
mem_array[6195] = 16'hd6e6;
mem_array[6194] = 16'h3e50;
mem_array[6197] = 16'hbf76;
mem_array[6196] = 16'hbde1;
mem_array[6199] = 16'h72ef;
mem_array[6198] = 16'hbee1;
mem_array[6201] = 16'h4fce;
mem_array[6200] = 16'hbd93;
mem_array[6203] = 16'hb240;
mem_array[6202] = 16'h3c96;
mem_array[6205] = 16'h4d3a;
mem_array[6204] = 16'hbe0c;
mem_array[6207] = 16'ha9b4;
mem_array[6206] = 16'hbea4;
mem_array[6209] = 16'h796f;
mem_array[6208] = 16'h3f3d;
mem_array[6211] = 16'h1743;
mem_array[6210] = 16'hbd43;
mem_array[6213] = 16'hb51f;
mem_array[6212] = 16'h3ed0;
mem_array[6215] = 16'hfda7;
mem_array[6214] = 16'h3df8;
mem_array[6217] = 16'h5489;
mem_array[6216] = 16'h3e92;
mem_array[6219] = 16'h29aa;
mem_array[6218] = 16'h3f2f;
mem_array[6221] = 16'h381f;
mem_array[6220] = 16'hbeef;
mem_array[6223] = 16'h4091;
mem_array[6222] = 16'h3d87;
mem_array[6225] = 16'h5f55;
mem_array[6224] = 16'h3e10;
mem_array[6227] = 16'h1535;
mem_array[6226] = 16'h3f55;
mem_array[6229] = 16'h5056;
mem_array[6228] = 16'hbed9;
mem_array[6231] = 16'h8993;
mem_array[6230] = 16'hbe1f;
mem_array[6233] = 16'h23f6;
mem_array[6232] = 16'hbee3;
mem_array[6235] = 16'he9d0;
mem_array[6234] = 16'h3efc;
mem_array[6237] = 16'ha178;
mem_array[6236] = 16'hbcc5;
mem_array[6239] = 16'hd6f3;
mem_array[6238] = 16'hbbfb;
mem_array[6241] = 16'h40ba;
mem_array[6240] = 16'h3eca;
mem_array[6243] = 16'h81e6;
mem_array[6242] = 16'hbe4b;
mem_array[6245] = 16'h865c;
mem_array[6244] = 16'hbf94;
mem_array[6247] = 16'h6398;
mem_array[6246] = 16'hbe5e;
mem_array[6249] = 16'h2da2;
mem_array[6248] = 16'h3eac;
mem_array[6251] = 16'h4078;
mem_array[6250] = 16'h3b94;
mem_array[6253] = 16'hb093;
mem_array[6252] = 16'h3eab;
mem_array[6255] = 16'h91db;
mem_array[6254] = 16'h3f8e;
mem_array[6257] = 16'hfe01;
mem_array[6256] = 16'hbeec;
mem_array[6259] = 16'h00ab;
mem_array[6258] = 16'hbf14;
mem_array[6261] = 16'h5cae;
mem_array[6260] = 16'hbcb0;
mem_array[6263] = 16'h7ff7;
mem_array[6262] = 16'h3db1;
mem_array[6265] = 16'h8f79;
mem_array[6264] = 16'hbec7;
mem_array[6267] = 16'h7634;
mem_array[6266] = 16'hbeff;
mem_array[6269] = 16'hbac0;
mem_array[6268] = 16'h3e36;
mem_array[6271] = 16'h627a;
mem_array[6270] = 16'hbdff;
mem_array[6273] = 16'hb784;
mem_array[6272] = 16'hbeaa;
mem_array[6275] = 16'h2fda;
mem_array[6274] = 16'hbdb4;
mem_array[6277] = 16'h7a6c;
mem_array[6276] = 16'h3ed0;
mem_array[6279] = 16'h1222;
mem_array[6278] = 16'h3e6a;
mem_array[6281] = 16'hebfe;
mem_array[6280] = 16'hbee5;
mem_array[6283] = 16'h198e;
mem_array[6282] = 16'h3ec5;
mem_array[6285] = 16'hf219;
mem_array[6284] = 16'h3c5e;
mem_array[6287] = 16'h9726;
mem_array[6286] = 16'h3d3b;
mem_array[6289] = 16'h90d0;
mem_array[6288] = 16'hbebf;
mem_array[6291] = 16'hf080;
mem_array[6290] = 16'h3b8c;
mem_array[6293] = 16'h281d;
mem_array[6292] = 16'h3e6a;
mem_array[6295] = 16'ha344;
mem_array[6294] = 16'h3f53;
mem_array[6297] = 16'h8460;
mem_array[6296] = 16'h3ec4;
mem_array[6299] = 16'h25ce;
mem_array[6298] = 16'hbf2c;
mem_array[6301] = 16'h81ac;
mem_array[6300] = 16'h3d9c;
mem_array[6303] = 16'h65a3;
mem_array[6302] = 16'hbe30;
mem_array[6305] = 16'h68e5;
mem_array[6304] = 16'hbf2b;
mem_array[6307] = 16'h1e75;
mem_array[6306] = 16'hbe63;
mem_array[6309] = 16'h4d71;
mem_array[6308] = 16'h3f57;
mem_array[6311] = 16'h456a;
mem_array[6310] = 16'h3e94;
mem_array[6313] = 16'ha9a2;
mem_array[6312] = 16'hbf95;
mem_array[6315] = 16'h66fe;
mem_array[6314] = 16'h3e88;
mem_array[6317] = 16'h231d;
mem_array[6316] = 16'h3d7f;
mem_array[6319] = 16'h9294;
mem_array[6318] = 16'hbf46;
mem_array[6321] = 16'h042f;
mem_array[6320] = 16'hbd10;
mem_array[6323] = 16'h1510;
mem_array[6322] = 16'h3ccf;
mem_array[6325] = 16'h4e81;
mem_array[6324] = 16'h3a9a;
mem_array[6327] = 16'h001f;
mem_array[6326] = 16'hbf2b;
mem_array[6329] = 16'hded2;
mem_array[6328] = 16'h3ef4;
mem_array[6331] = 16'hc51e;
mem_array[6330] = 16'hbae7;
mem_array[6333] = 16'h3719;
mem_array[6332] = 16'hbef5;
mem_array[6335] = 16'h1980;
mem_array[6334] = 16'h3ee7;
mem_array[6337] = 16'hc650;
mem_array[6336] = 16'hbf02;
mem_array[6339] = 16'h2ee7;
mem_array[6338] = 16'h3ecf;
mem_array[6341] = 16'h5fc8;
mem_array[6340] = 16'h3f32;
mem_array[6343] = 16'h2ee1;
mem_array[6342] = 16'h3f23;
mem_array[6345] = 16'hd8dd;
mem_array[6344] = 16'h3e03;
mem_array[6347] = 16'hf782;
mem_array[6346] = 16'h3ef7;
mem_array[6349] = 16'hb84c;
mem_array[6348] = 16'h3d19;
mem_array[6351] = 16'h9392;
mem_array[6350] = 16'hbd51;
mem_array[6353] = 16'hba0f;
mem_array[6352] = 16'h3d31;
mem_array[6355] = 16'hdc92;
mem_array[6354] = 16'h3ebd;
mem_array[6357] = 16'h6ed7;
mem_array[6356] = 16'h3e43;
mem_array[6359] = 16'h453c;
mem_array[6358] = 16'hbf07;
mem_array[6361] = 16'hbfeb;
mem_array[6360] = 16'h3eca;
mem_array[6363] = 16'h60fd;
mem_array[6362] = 16'h3d07;
mem_array[6365] = 16'h8b11;
mem_array[6364] = 16'h3d7a;
mem_array[6367] = 16'hfe94;
mem_array[6366] = 16'hbf26;
mem_array[6369] = 16'h3cee;
mem_array[6368] = 16'h3f42;
mem_array[6371] = 16'h65c7;
mem_array[6370] = 16'h3da2;
mem_array[6373] = 16'ha922;
mem_array[6372] = 16'hbfa5;
mem_array[6375] = 16'h8b7e;
mem_array[6374] = 16'hbe8d;
mem_array[6377] = 16'he00f;
mem_array[6376] = 16'hbdac;
mem_array[6379] = 16'hdcea;
mem_array[6378] = 16'h3f8f;
mem_array[6381] = 16'h7271;
mem_array[6380] = 16'hbdd8;
mem_array[6383] = 16'hfe38;
mem_array[6382] = 16'hbc26;
mem_array[6385] = 16'h8f61;
mem_array[6384] = 16'hbe88;
mem_array[6387] = 16'hb247;
mem_array[6386] = 16'h3f2c;
mem_array[6389] = 16'h3cc8;
mem_array[6388] = 16'hbdba;
mem_array[6391] = 16'h4069;
mem_array[6390] = 16'h3cf4;
mem_array[6393] = 16'h46d4;
mem_array[6392] = 16'h3f30;
mem_array[6395] = 16'h928c;
mem_array[6394] = 16'h3eeb;
mem_array[6397] = 16'hbfba;
mem_array[6396] = 16'hbfb3;
mem_array[6399] = 16'h744b;
mem_array[6398] = 16'h3efe;
mem_array[6401] = 16'h45f2;
mem_array[6400] = 16'hbd18;
mem_array[6403] = 16'ha8c6;
mem_array[6402] = 16'h3d0e;
mem_array[6405] = 16'h2921;
mem_array[6404] = 16'h3ec0;
mem_array[6407] = 16'hcdb9;
mem_array[6406] = 16'h3eb0;
mem_array[6409] = 16'h58fb;
mem_array[6408] = 16'h3eb5;
mem_array[6411] = 16'h894f;
mem_array[6410] = 16'h3e71;
mem_array[6413] = 16'hc475;
mem_array[6412] = 16'h3ec5;
mem_array[6415] = 16'h7cd7;
mem_array[6414] = 16'h3c5d;
mem_array[6417] = 16'h9e3c;
mem_array[6416] = 16'h3d8d;
mem_array[6419] = 16'hd8d4;
mem_array[6418] = 16'hbd85;
mem_array[6421] = 16'hc972;
mem_array[6420] = 16'h3eac;
mem_array[6423] = 16'h57f3;
mem_array[6422] = 16'h3ee6;
mem_array[6425] = 16'hcc76;
mem_array[6424] = 16'h3f72;
mem_array[6427] = 16'hacf2;
mem_array[6426] = 16'hbe32;
mem_array[6429] = 16'h328a;
mem_array[6428] = 16'h3f03;
mem_array[6431] = 16'hee65;
mem_array[6430] = 16'hbe02;
mem_array[6433] = 16'hbb78;
mem_array[6432] = 16'hbfcf;
mem_array[6435] = 16'hbebe;
mem_array[6434] = 16'h3f28;
mem_array[6437] = 16'he45f;
mem_array[6436] = 16'h3def;
mem_array[6439] = 16'ha154;
mem_array[6438] = 16'h3c7f;
mem_array[6441] = 16'h417e;
mem_array[6440] = 16'h3dd2;
mem_array[6443] = 16'h5b69;
mem_array[6442] = 16'hbd88;
mem_array[6445] = 16'hd0e5;
mem_array[6444] = 16'hbeb3;
mem_array[6447] = 16'h379d;
mem_array[6446] = 16'hbf08;
mem_array[6449] = 16'h8ee2;
mem_array[6448] = 16'hbea7;
mem_array[6451] = 16'h645d;
mem_array[6450] = 16'h3e97;
mem_array[6453] = 16'h203c;
mem_array[6452] = 16'h3eb9;
mem_array[6455] = 16'h1855;
mem_array[6454] = 16'h3e5a;
mem_array[6457] = 16'h2f8f;
mem_array[6456] = 16'hbcf4;
mem_array[6459] = 16'hf489;
mem_array[6458] = 16'hbebb;
mem_array[6461] = 16'h92e7;
mem_array[6460] = 16'hbe95;
mem_array[6463] = 16'hf0d0;
mem_array[6462] = 16'hbd5e;
mem_array[6465] = 16'hba14;
mem_array[6464] = 16'hbf96;
mem_array[6467] = 16'hfbf6;
mem_array[6466] = 16'h3f75;
mem_array[6469] = 16'h3edd;
mem_array[6468] = 16'hbf13;
mem_array[6471] = 16'hd19e;
mem_array[6470] = 16'h3c51;
mem_array[6473] = 16'h93ee;
mem_array[6472] = 16'h3d37;
mem_array[6475] = 16'h1e29;
mem_array[6474] = 16'h3d03;
mem_array[6477] = 16'hfde3;
mem_array[6476] = 16'h3d4d;
mem_array[6479] = 16'h20f4;
mem_array[6478] = 16'h3e67;
mem_array[6481] = 16'he1cb;
mem_array[6480] = 16'hbeb4;
mem_array[6483] = 16'h2758;
mem_array[6482] = 16'h3ebb;
mem_array[6485] = 16'h43e6;
mem_array[6484] = 16'hbd10;
mem_array[6487] = 16'h6b40;
mem_array[6486] = 16'hbe06;
mem_array[6489] = 16'hda47;
mem_array[6488] = 16'h3e5c;
mem_array[6491] = 16'h090e;
mem_array[6490] = 16'h3eca;
mem_array[6493] = 16'h9ca0;
mem_array[6492] = 16'hbf07;
mem_array[6495] = 16'h9974;
mem_array[6494] = 16'h3ea3;
mem_array[6497] = 16'he517;
mem_array[6496] = 16'h3ed8;
mem_array[6499] = 16'h0f91;
mem_array[6498] = 16'hbd99;
mem_array[6501] = 16'h2949;
mem_array[6500] = 16'hbcb1;
mem_array[6503] = 16'h71a3;
mem_array[6502] = 16'hbc08;
mem_array[6505] = 16'h29c4;
mem_array[6504] = 16'hbf09;
mem_array[6507] = 16'h5e45;
mem_array[6506] = 16'hbde6;
mem_array[6509] = 16'h6ebb;
mem_array[6508] = 16'hbf1a;
mem_array[6511] = 16'h5582;
mem_array[6510] = 16'h3e6e;
mem_array[6513] = 16'hd93d;
mem_array[6512] = 16'hbe58;
mem_array[6515] = 16'h2c18;
mem_array[6514] = 16'h3edc;
mem_array[6517] = 16'h7769;
mem_array[6516] = 16'h3d5c;
mem_array[6519] = 16'h43b6;
mem_array[6518] = 16'h3dcc;
mem_array[6521] = 16'h6b1e;
mem_array[6520] = 16'hbea2;
mem_array[6523] = 16'hb5a2;
mem_array[6522] = 16'h3f21;
mem_array[6525] = 16'h5dbd;
mem_array[6524] = 16'hbf68;
mem_array[6527] = 16'h717a;
mem_array[6526] = 16'h3d30;
mem_array[6529] = 16'hfc3d;
mem_array[6528] = 16'hbe83;
mem_array[6531] = 16'hf95a;
mem_array[6530] = 16'h3d8d;
mem_array[6533] = 16'h3b8e;
mem_array[6532] = 16'h3e87;
mem_array[6535] = 16'hbea0;
mem_array[6534] = 16'hbd29;
mem_array[6537] = 16'h03e6;
mem_array[6536] = 16'h3e81;
mem_array[6539] = 16'hd91b;
mem_array[6538] = 16'hbf00;
mem_array[6541] = 16'h8220;
mem_array[6540] = 16'hbeac;
mem_array[6543] = 16'hb51b;
mem_array[6542] = 16'h3d8b;
mem_array[6545] = 16'h9c67;
mem_array[6544] = 16'hbbd3;
mem_array[6547] = 16'hcec1;
mem_array[6546] = 16'h3ebb;
mem_array[6549] = 16'h47ef;
mem_array[6548] = 16'h3d19;
mem_array[6551] = 16'h9cd7;
mem_array[6550] = 16'hbebc;
mem_array[6553] = 16'hc499;
mem_array[6552] = 16'h3e6b;
mem_array[6555] = 16'h9fd0;
mem_array[6554] = 16'h3ebf;
mem_array[6557] = 16'h7936;
mem_array[6556] = 16'h3f22;
mem_array[6559] = 16'h8f9a;
mem_array[6558] = 16'hbdc2;
mem_array[6561] = 16'h8a2f;
mem_array[6560] = 16'hbd93;
mem_array[6563] = 16'he406;
mem_array[6562] = 16'h3d49;
mem_array[6565] = 16'h04f7;
mem_array[6564] = 16'hbd8b;
mem_array[6567] = 16'haad8;
mem_array[6566] = 16'h3f1b;
mem_array[6569] = 16'h4fb5;
mem_array[6568] = 16'h3de3;
mem_array[6571] = 16'h8cd8;
mem_array[6570] = 16'h3e10;
mem_array[6573] = 16'h7751;
mem_array[6572] = 16'hbddb;
mem_array[6575] = 16'h65d8;
mem_array[6574] = 16'h3e21;
mem_array[6577] = 16'h28c2;
mem_array[6576] = 16'h3dcf;
mem_array[6579] = 16'hd550;
mem_array[6578] = 16'h39e9;
mem_array[6581] = 16'hf453;
mem_array[6580] = 16'h3db4;
mem_array[6583] = 16'h3218;
mem_array[6582] = 16'hbef1;
mem_array[6585] = 16'h837e;
mem_array[6584] = 16'hbeb2;
mem_array[6587] = 16'h8f7a;
mem_array[6586] = 16'hbe35;
mem_array[6589] = 16'ha56a;
mem_array[6588] = 16'h3db5;
mem_array[6591] = 16'h41db;
mem_array[6590] = 16'h3c61;
mem_array[6593] = 16'h914b;
mem_array[6592] = 16'h3d9d;
mem_array[6595] = 16'hb28c;
mem_array[6594] = 16'hbefd;
mem_array[6597] = 16'h856b;
mem_array[6596] = 16'h3ef9;
mem_array[6599] = 16'h81a5;
mem_array[6598] = 16'h3e91;
mem_array[6601] = 16'h023a;
mem_array[6600] = 16'hbe30;
mem_array[6603] = 16'hbbbe;
mem_array[6602] = 16'hbd01;
mem_array[6605] = 16'hb6b9;
mem_array[6604] = 16'h3dc7;
mem_array[6607] = 16'hbc24;
mem_array[6606] = 16'hbcf1;
mem_array[6609] = 16'hc2e2;
mem_array[6608] = 16'h3cf7;
mem_array[6611] = 16'h8c5e;
mem_array[6610] = 16'hbd78;
mem_array[6613] = 16'hdc44;
mem_array[6612] = 16'hbd69;
mem_array[6615] = 16'h067e;
mem_array[6614] = 16'hbdd7;
mem_array[6617] = 16'hb3d0;
mem_array[6616] = 16'h3d0f;
mem_array[6619] = 16'h4c27;
mem_array[6618] = 16'hbd98;
mem_array[6621] = 16'hbdf6;
mem_array[6620] = 16'hbd7e;
mem_array[6623] = 16'h062f;
mem_array[6622] = 16'hbc18;
mem_array[6625] = 16'hd443;
mem_array[6624] = 16'h3e67;
mem_array[6627] = 16'h07db;
mem_array[6626] = 16'hbdce;
mem_array[6629] = 16'hcab4;
mem_array[6628] = 16'hbcaa;
mem_array[6631] = 16'hec8e;
mem_array[6630] = 16'hbe84;
mem_array[6633] = 16'h0351;
mem_array[6632] = 16'h3d05;
mem_array[6635] = 16'hf3b4;
mem_array[6634] = 16'hbc30;
mem_array[6637] = 16'h13c5;
mem_array[6636] = 16'hbc08;
mem_array[6639] = 16'h6bf0;
mem_array[6638] = 16'h3d28;
mem_array[6641] = 16'h3f0c;
mem_array[6640] = 16'hbd98;
mem_array[6643] = 16'h68b8;
mem_array[6642] = 16'h3e6b;
mem_array[6645] = 16'h9363;
mem_array[6644] = 16'h3d23;
mem_array[6647] = 16'h1240;
mem_array[6646] = 16'h3edd;
mem_array[6649] = 16'h50dd;
mem_array[6648] = 16'hbdbb;
mem_array[6651] = 16'h42d2;
mem_array[6650] = 16'h3d12;
mem_array[6653] = 16'hd58c;
mem_array[6652] = 16'hbe92;
mem_array[6655] = 16'h46a0;
mem_array[6654] = 16'h3c63;
mem_array[6657] = 16'habdc;
mem_array[6656] = 16'hbdcc;
mem_array[6659] = 16'hc64b;
mem_array[6658] = 16'h3e93;
mem_array[6661] = 16'h5811;
mem_array[6660] = 16'h3d6b;
mem_array[6663] = 16'had57;
mem_array[6662] = 16'hbd57;
mem_array[6665] = 16'h8091;
mem_array[6664] = 16'h3c58;
mem_array[6667] = 16'h4750;
mem_array[6666] = 16'h3d2c;
mem_array[6669] = 16'h3b2b;
mem_array[6668] = 16'hbd4e;
mem_array[6671] = 16'h9125;
mem_array[6670] = 16'hbc16;
mem_array[6673] = 16'h8f00;
mem_array[6672] = 16'hbce6;
mem_array[6675] = 16'h4b62;
mem_array[6674] = 16'hbca7;
mem_array[6677] = 16'h5e2b;
mem_array[6676] = 16'hbd1b;
mem_array[6679] = 16'h9dda;
mem_array[6678] = 16'hbd7d;
mem_array[6681] = 16'h7d31;
mem_array[6680] = 16'hbc94;
mem_array[6683] = 16'h1c70;
mem_array[6682] = 16'h3ae2;
mem_array[6685] = 16'h7117;
mem_array[6684] = 16'hbce1;
mem_array[6687] = 16'h3b26;
mem_array[6686] = 16'hbdc1;
mem_array[6689] = 16'h705d;
mem_array[6688] = 16'h3c1b;
mem_array[6691] = 16'h7f11;
mem_array[6690] = 16'h3bc4;
mem_array[6693] = 16'h3135;
mem_array[6692] = 16'hbc96;
mem_array[6695] = 16'h50b4;
mem_array[6694] = 16'h3c20;
mem_array[6697] = 16'h97e3;
mem_array[6696] = 16'h3cdb;
mem_array[6699] = 16'ha4fb;
mem_array[6698] = 16'h3dc6;
mem_array[6701] = 16'h9d33;
mem_array[6700] = 16'hbd0e;
mem_array[6703] = 16'h4ab3;
mem_array[6702] = 16'h3d26;
mem_array[6705] = 16'ha016;
mem_array[6704] = 16'h3d52;
mem_array[6707] = 16'h7d2a;
mem_array[6706] = 16'hbca4;
mem_array[6709] = 16'h3548;
mem_array[6708] = 16'h3d50;
mem_array[6711] = 16'h37d3;
mem_array[6710] = 16'h3bea;
mem_array[6713] = 16'hf99c;
mem_array[6712] = 16'hbb2b;
mem_array[6715] = 16'h237d;
mem_array[6714] = 16'h3ce7;
mem_array[6717] = 16'h2a67;
mem_array[6716] = 16'hbc84;
mem_array[6719] = 16'h426d;
mem_array[6718] = 16'hbcef;
mem_array[6721] = 16'hc25d;
mem_array[6720] = 16'hbdcf;
mem_array[6723] = 16'hfd53;
mem_array[6722] = 16'hbc73;
mem_array[6725] = 16'heeef;
mem_array[6724] = 16'hbd8c;
mem_array[6727] = 16'h17e1;
mem_array[6726] = 16'h3ccc;
mem_array[6729] = 16'hd488;
mem_array[6728] = 16'hbd32;
mem_array[6731] = 16'h90f7;
mem_array[6730] = 16'h3d78;
mem_array[6733] = 16'h1905;
mem_array[6732] = 16'hbbd3;
mem_array[6735] = 16'h501f;
mem_array[6734] = 16'h3d8c;
mem_array[6737] = 16'h3ba3;
mem_array[6736] = 16'h3c61;
mem_array[6739] = 16'h6bfa;
mem_array[6738] = 16'hbc62;
mem_array[6741] = 16'h7c9d;
mem_array[6740] = 16'h3d9c;
mem_array[6743] = 16'h4f90;
mem_array[6742] = 16'h3cc2;
mem_array[6745] = 16'h148c;
mem_array[6744] = 16'h3d5d;
mem_array[6747] = 16'h4259;
mem_array[6746] = 16'hbdd7;
mem_array[6749] = 16'h6fe5;
mem_array[6748] = 16'h3d24;
mem_array[6751] = 16'h3d5b;
mem_array[6750] = 16'hbca1;
mem_array[6753] = 16'h8f27;
mem_array[6752] = 16'hbd11;
mem_array[6755] = 16'hfbe0;
mem_array[6754] = 16'hbd04;
mem_array[6757] = 16'hd15d;
mem_array[6756] = 16'hbcac;
mem_array[6759] = 16'hfa09;
mem_array[6758] = 16'hbc31;
mem_array[6761] = 16'hec8c;
mem_array[6760] = 16'h3d81;
mem_array[6763] = 16'hbc88;
mem_array[6762] = 16'h3d74;
mem_array[6765] = 16'h9ed3;
mem_array[6764] = 16'hbcfc;
mem_array[6767] = 16'h30e2;
mem_array[6766] = 16'h3ba2;
mem_array[6769] = 16'hd4aa;
mem_array[6768] = 16'h3c0e;
mem_array[6771] = 16'hb3c8;
mem_array[6770] = 16'h3d0c;
mem_array[6773] = 16'hf0ce;
mem_array[6772] = 16'hbbc3;
mem_array[6775] = 16'h1002;
mem_array[6774] = 16'h3dca;
mem_array[6777] = 16'h1f6f;
mem_array[6776] = 16'hbd9b;
mem_array[6779] = 16'ha24a;
mem_array[6778] = 16'h3d28;
mem_array[6781] = 16'h3252;
mem_array[6780] = 16'h3d00;
mem_array[6783] = 16'haeac;
mem_array[6782] = 16'hbb71;
mem_array[6785] = 16'h8b8b;
mem_array[6784] = 16'h3b88;
mem_array[6787] = 16'hd13c;
mem_array[6786] = 16'hbd15;
mem_array[6789] = 16'hef79;
mem_array[6788] = 16'hbd4b;
mem_array[6791] = 16'h8760;
mem_array[6790] = 16'h3d41;
mem_array[6793] = 16'hbf1a;
mem_array[6792] = 16'hbec3;
mem_array[6795] = 16'h0f70;
mem_array[6794] = 16'hbd3a;
mem_array[6797] = 16'h77a0;
mem_array[6796] = 16'h3d71;
mem_array[6799] = 16'h325a;
mem_array[6798] = 16'hbd04;
mem_array[6801] = 16'h9bea;
mem_array[6800] = 16'h3d19;
mem_array[6803] = 16'h4c09;
mem_array[6802] = 16'hbd81;
mem_array[6805] = 16'heb89;
mem_array[6804] = 16'h3bf1;
mem_array[6807] = 16'ha0ab;
mem_array[6806] = 16'hbd89;
mem_array[6809] = 16'hbca6;
mem_array[6808] = 16'hbcb3;
mem_array[6811] = 16'h98d9;
mem_array[6810] = 16'hbea7;
mem_array[6813] = 16'h51d6;
mem_array[6812] = 16'hbdb7;
mem_array[6815] = 16'haa27;
mem_array[6814] = 16'h3d7b;
mem_array[6817] = 16'hb0bf;
mem_array[6816] = 16'hbbd6;
mem_array[6819] = 16'h6ecc;
mem_array[6818] = 16'hbadc;
mem_array[6821] = 16'h8f6b;
mem_array[6820] = 16'h3c10;
mem_array[6823] = 16'h4eff;
mem_array[6822] = 16'hbe2a;
mem_array[6825] = 16'he9b2;
mem_array[6824] = 16'h3cf8;
mem_array[6827] = 16'h4116;
mem_array[6826] = 16'h3ee4;
mem_array[6829] = 16'hceb5;
mem_array[6828] = 16'hbf0e;
mem_array[6831] = 16'h4c3f;
mem_array[6830] = 16'h3d8a;
mem_array[6833] = 16'h5f3c;
mem_array[6832] = 16'hbf04;
mem_array[6835] = 16'hb459;
mem_array[6834] = 16'hbcb9;
mem_array[6837] = 16'h05fc;
mem_array[6836] = 16'hbe29;
mem_array[6839] = 16'hde07;
mem_array[6838] = 16'h3e01;
mem_array[6841] = 16'h8180;
mem_array[6840] = 16'h3ed8;
mem_array[6843] = 16'h3fc2;
mem_array[6842] = 16'h3dc6;
mem_array[6845] = 16'h49b5;
mem_array[6844] = 16'h3df6;
mem_array[6847] = 16'h9618;
mem_array[6846] = 16'h3d18;
mem_array[6849] = 16'h69f5;
mem_array[6848] = 16'h3d34;
mem_array[6851] = 16'h2d62;
mem_array[6850] = 16'h3d8d;
mem_array[6853] = 16'h288d;
mem_array[6852] = 16'h3e50;
mem_array[6855] = 16'h9cb2;
mem_array[6854] = 16'h3e88;
mem_array[6857] = 16'ha96a;
mem_array[6856] = 16'h3cdd;
mem_array[6859] = 16'h5336;
mem_array[6858] = 16'h3f38;
mem_array[6861] = 16'h7dd3;
mem_array[6860] = 16'h3c6c;
mem_array[6863] = 16'h9767;
mem_array[6862] = 16'hba3e;
mem_array[6865] = 16'h02e1;
mem_array[6864] = 16'hbe0d;
mem_array[6867] = 16'h05ad;
mem_array[6866] = 16'h3e2e;
mem_array[6869] = 16'hac8b;
mem_array[6868] = 16'hbd33;
mem_array[6871] = 16'hd7d9;
mem_array[6870] = 16'h3f51;
mem_array[6873] = 16'h9aa7;
mem_array[6872] = 16'hbcce;
mem_array[6875] = 16'ha00f;
mem_array[6874] = 16'hbc6f;
mem_array[6877] = 16'h2b49;
mem_array[6876] = 16'h3c7b;
mem_array[6879] = 16'h7320;
mem_array[6878] = 16'hbc17;
mem_array[6881] = 16'h3a05;
mem_array[6880] = 16'hbe66;
mem_array[6883] = 16'hce3d;
mem_array[6882] = 16'hbf33;
mem_array[6885] = 16'h6f0d;
mem_array[6884] = 16'hbf2d;
mem_array[6887] = 16'h8dca;
mem_array[6886] = 16'hbf82;
mem_array[6889] = 16'h5fc9;
mem_array[6888] = 16'h3d49;
mem_array[6891] = 16'haf2e;
mem_array[6890] = 16'h3d4f;
mem_array[6893] = 16'habda;
mem_array[6892] = 16'h3e4e;
mem_array[6895] = 16'h2299;
mem_array[6894] = 16'hbd67;
mem_array[6897] = 16'hb5a3;
mem_array[6896] = 16'h3da5;
mem_array[6899] = 16'h2001;
mem_array[6898] = 16'hbeaf;
mem_array[6901] = 16'he0c8;
mem_array[6900] = 16'h3ec7;
mem_array[6903] = 16'h7bda;
mem_array[6902] = 16'hbce5;
mem_array[6905] = 16'hfa94;
mem_array[6904] = 16'hbeae;
mem_array[6907] = 16'hcd6e;
mem_array[6906] = 16'h3e59;
mem_array[6909] = 16'h9652;
mem_array[6908] = 16'hbe02;
mem_array[6911] = 16'h99ed;
mem_array[6910] = 16'h3cd4;
mem_array[6913] = 16'hf4bb;
mem_array[6912] = 16'hbe6b;
mem_array[6915] = 16'ha42c;
mem_array[6914] = 16'h3f48;
mem_array[6917] = 16'h12ef;
mem_array[6916] = 16'hbd9e;
mem_array[6919] = 16'h123d;
mem_array[6918] = 16'h3f38;
mem_array[6921] = 16'hc929;
mem_array[6920] = 16'hbd6f;
mem_array[6923] = 16'h7886;
mem_array[6922] = 16'hbd2b;
mem_array[6925] = 16'had4e;
mem_array[6924] = 16'h3c88;
mem_array[6927] = 16'h2754;
mem_array[6926] = 16'hbeac;
mem_array[6929] = 16'he28e;
mem_array[6928] = 16'h3e12;
mem_array[6931] = 16'ha534;
mem_array[6930] = 16'h3f26;
mem_array[6933] = 16'hd3df;
mem_array[6932] = 16'hbd87;
mem_array[6935] = 16'hb162;
mem_array[6934] = 16'hbf09;
mem_array[6937] = 16'hdffc;
mem_array[6936] = 16'h3e83;
mem_array[6939] = 16'h05a3;
mem_array[6938] = 16'hbe8f;
mem_array[6941] = 16'h5b01;
mem_array[6940] = 16'hbdab;
mem_array[6943] = 16'h9573;
mem_array[6942] = 16'h3f20;
mem_array[6945] = 16'h3092;
mem_array[6944] = 16'hbf29;
mem_array[6947] = 16'h0450;
mem_array[6946] = 16'h3ad8;
mem_array[6949] = 16'h566e;
mem_array[6948] = 16'hbf04;
mem_array[6951] = 16'hd5f1;
mem_array[6950] = 16'h3e9f;
mem_array[6953] = 16'h6b05;
mem_array[6952] = 16'h3e08;
mem_array[6955] = 16'hcd0c;
mem_array[6954] = 16'h3e9f;
mem_array[6957] = 16'h9e1b;
mem_array[6956] = 16'h3e19;
mem_array[6959] = 16'hf0b2;
mem_array[6958] = 16'hbf80;
mem_array[6961] = 16'ha266;
mem_array[6960] = 16'hbe88;
mem_array[6963] = 16'h0c38;
mem_array[6962] = 16'hbead;
mem_array[6965] = 16'h6b38;
mem_array[6964] = 16'h3e38;
mem_array[6967] = 16'hdce3;
mem_array[6966] = 16'h3ec6;
mem_array[6969] = 16'hbbc3;
mem_array[6968] = 16'h3f10;
mem_array[6971] = 16'h4e8d;
mem_array[6970] = 16'hbeba;
mem_array[6973] = 16'h9665;
mem_array[6972] = 16'h3f49;
mem_array[6975] = 16'h04ea;
mem_array[6974] = 16'h3e3d;
mem_array[6977] = 16'hadb4;
mem_array[6976] = 16'h3e9f;
mem_array[6979] = 16'ha8bc;
mem_array[6978] = 16'hbcde;
mem_array[6981] = 16'hc810;
mem_array[6980] = 16'h3bb3;
mem_array[6983] = 16'h25eb;
mem_array[6982] = 16'hbc93;
mem_array[6985] = 16'ha39d;
mem_array[6984] = 16'hbf9f;
mem_array[6987] = 16'h95dd;
mem_array[6986] = 16'h3e48;
mem_array[6989] = 16'hecfb;
mem_array[6988] = 16'h3f17;
mem_array[6991] = 16'h9c42;
mem_array[6990] = 16'hbe8f;
mem_array[6993] = 16'h7164;
mem_array[6992] = 16'h3ec7;
mem_array[6995] = 16'h77a7;
mem_array[6994] = 16'hbe32;
mem_array[6997] = 16'hb15f;
mem_array[6996] = 16'hbf0f;
mem_array[6999] = 16'h23fb;
mem_array[6998] = 16'h3e1f;
mem_array[7001] = 16'h5912;
mem_array[7000] = 16'h3e1d;
mem_array[7003] = 16'h6b57;
mem_array[7002] = 16'h3edb;
mem_array[7005] = 16'hfe77;
mem_array[7004] = 16'h3c88;
mem_array[7007] = 16'h488f;
mem_array[7006] = 16'h3f1b;
mem_array[7009] = 16'h2c54;
mem_array[7008] = 16'hbdb0;
mem_array[7011] = 16'h7620;
mem_array[7010] = 16'h3e12;
mem_array[7013] = 16'hec14;
mem_array[7012] = 16'h3f22;
mem_array[7015] = 16'heaca;
mem_array[7014] = 16'h3f39;
mem_array[7017] = 16'hfb55;
mem_array[7016] = 16'h3e94;
mem_array[7019] = 16'h0726;
mem_array[7018] = 16'h3df4;
mem_array[7021] = 16'h6096;
mem_array[7020] = 16'hbe83;
mem_array[7023] = 16'h5406;
mem_array[7022] = 16'h3dec;
mem_array[7025] = 16'h366d;
mem_array[7024] = 16'h3dc8;
mem_array[7027] = 16'hd19d;
mem_array[7026] = 16'hbf28;
mem_array[7029] = 16'hb496;
mem_array[7028] = 16'h3f0f;
mem_array[7031] = 16'hd854;
mem_array[7030] = 16'hbf19;
mem_array[7033] = 16'hbc3f;
mem_array[7032] = 16'h3fa8;
mem_array[7035] = 16'hb817;
mem_array[7034] = 16'h3e9e;
mem_array[7037] = 16'h2d0c;
mem_array[7036] = 16'h3dfd;
mem_array[7039] = 16'hc845;
mem_array[7038] = 16'h3f32;
mem_array[7041] = 16'h5cc7;
mem_array[7040] = 16'hbc51;
mem_array[7043] = 16'h10de;
mem_array[7042] = 16'h3d10;
mem_array[7045] = 16'h03d7;
mem_array[7044] = 16'hbf89;
mem_array[7047] = 16'h40bc;
mem_array[7046] = 16'hbefb;
mem_array[7049] = 16'hcdb0;
mem_array[7048] = 16'h3f33;
mem_array[7051] = 16'h31e0;
mem_array[7050] = 16'h3e1c;
mem_array[7053] = 16'h0e18;
mem_array[7052] = 16'h3f16;
mem_array[7055] = 16'h7a33;
mem_array[7054] = 16'h3f3d;
mem_array[7057] = 16'hc3b4;
mem_array[7056] = 16'hbcb3;
mem_array[7059] = 16'h4ab0;
mem_array[7058] = 16'h3f43;
mem_array[7061] = 16'h5cbd;
mem_array[7060] = 16'h3f13;
mem_array[7063] = 16'h7985;
mem_array[7062] = 16'hbe7c;
mem_array[7065] = 16'h9f57;
mem_array[7064] = 16'hbe55;
mem_array[7067] = 16'h9670;
mem_array[7066] = 16'hbf40;
mem_array[7069] = 16'hb598;
mem_array[7068] = 16'h3f62;
mem_array[7071] = 16'h0cc3;
mem_array[7070] = 16'h3f1d;
mem_array[7073] = 16'h0bf6;
mem_array[7072] = 16'h3efe;
mem_array[7075] = 16'h4793;
mem_array[7074] = 16'h3f56;
mem_array[7077] = 16'h34c2;
mem_array[7076] = 16'h3dcc;
mem_array[7079] = 16'h89f2;
mem_array[7078] = 16'hbe8a;
mem_array[7081] = 16'h1094;
mem_array[7080] = 16'hbe41;
mem_array[7083] = 16'h9f44;
mem_array[7082] = 16'h3ec6;
mem_array[7085] = 16'h84e8;
mem_array[7084] = 16'h3eb8;
mem_array[7087] = 16'h6ca4;
mem_array[7086] = 16'hbf33;
mem_array[7089] = 16'hb8bf;
mem_array[7088] = 16'h3f03;
mem_array[7091] = 16'hc270;
mem_array[7090] = 16'hbf88;
mem_array[7093] = 16'h9c52;
mem_array[7092] = 16'h3f35;
mem_array[7095] = 16'h87ad;
mem_array[7094] = 16'h3ea5;
mem_array[7097] = 16'h62e0;
mem_array[7096] = 16'h3f1f;
mem_array[7099] = 16'h47fc;
mem_array[7098] = 16'hbe36;
mem_array[7101] = 16'he391;
mem_array[7100] = 16'h3b8d;
mem_array[7103] = 16'h6a61;
mem_array[7102] = 16'hbc0f;
mem_array[7105] = 16'h825f;
mem_array[7104] = 16'h3d71;
mem_array[7107] = 16'h1199;
mem_array[7106] = 16'h3e61;
mem_array[7109] = 16'h4012;
mem_array[7108] = 16'h3eb0;
mem_array[7111] = 16'hb262;
mem_array[7110] = 16'hbf09;
mem_array[7113] = 16'h5252;
mem_array[7112] = 16'hbc99;
mem_array[7115] = 16'he7be;
mem_array[7114] = 16'h3e68;
mem_array[7117] = 16'hee9a;
mem_array[7116] = 16'h3d80;
mem_array[7119] = 16'h6e06;
mem_array[7118] = 16'h3e32;
mem_array[7121] = 16'h801d;
mem_array[7120] = 16'h3e85;
mem_array[7123] = 16'h4abe;
mem_array[7122] = 16'h3e74;
mem_array[7125] = 16'h99e8;
mem_array[7124] = 16'hbee4;
mem_array[7127] = 16'h8c98;
mem_array[7126] = 16'hbe88;
mem_array[7129] = 16'h4877;
mem_array[7128] = 16'h3f0c;
mem_array[7131] = 16'hecd7;
mem_array[7130] = 16'h3f3d;
mem_array[7133] = 16'h3b7c;
mem_array[7132] = 16'h3d62;
mem_array[7135] = 16'heafb;
mem_array[7134] = 16'h3f34;
mem_array[7137] = 16'hec3f;
mem_array[7136] = 16'h3cad;
mem_array[7139] = 16'hfb10;
mem_array[7138] = 16'hbf88;
mem_array[7141] = 16'h6a9e;
mem_array[7140] = 16'h3f3a;
mem_array[7143] = 16'hd6d6;
mem_array[7142] = 16'hbf93;
mem_array[7145] = 16'h618e;
mem_array[7144] = 16'h3f20;
mem_array[7147] = 16'h663c;
mem_array[7146] = 16'hbee8;
mem_array[7149] = 16'h7a26;
mem_array[7148] = 16'h3f23;
mem_array[7151] = 16'h021a;
mem_array[7150] = 16'hbfab;
mem_array[7153] = 16'h4719;
mem_array[7152] = 16'h3cae;
mem_array[7155] = 16'hf939;
mem_array[7154] = 16'hbe0b;
mem_array[7157] = 16'h4e4c;
mem_array[7156] = 16'h3e68;
mem_array[7159] = 16'h04a8;
mem_array[7158] = 16'h3f18;
mem_array[7161] = 16'hd079;
mem_array[7160] = 16'h3d09;
mem_array[7163] = 16'hc4a3;
mem_array[7162] = 16'hbd54;
mem_array[7165] = 16'h4588;
mem_array[7164] = 16'h3dbc;
mem_array[7167] = 16'ha258;
mem_array[7166] = 16'h3f06;
mem_array[7169] = 16'hb197;
mem_array[7168] = 16'h3ea3;
mem_array[7171] = 16'hb001;
mem_array[7170] = 16'hbca7;
mem_array[7173] = 16'hef27;
mem_array[7172] = 16'h3f3b;
mem_array[7175] = 16'ha1a2;
mem_array[7174] = 16'h3f56;
mem_array[7177] = 16'h19bf;
mem_array[7176] = 16'hbdd3;
mem_array[7179] = 16'h3d6a;
mem_array[7178] = 16'h3e39;
mem_array[7181] = 16'ha5d5;
mem_array[7180] = 16'h3f0f;
mem_array[7183] = 16'h3adc;
mem_array[7182] = 16'h3f00;
mem_array[7185] = 16'h7230;
mem_array[7184] = 16'hbfb8;
mem_array[7187] = 16'h7179;
mem_array[7186] = 16'hbea8;
mem_array[7189] = 16'h5883;
mem_array[7188] = 16'h3f13;
mem_array[7191] = 16'h5775;
mem_array[7190] = 16'hbf07;
mem_array[7193] = 16'hc547;
mem_array[7192] = 16'hbcc5;
mem_array[7195] = 16'h493b;
mem_array[7194] = 16'h3eb4;
mem_array[7197] = 16'hf861;
mem_array[7196] = 16'hbe5e;
mem_array[7199] = 16'h266c;
mem_array[7198] = 16'hbf25;
mem_array[7201] = 16'hc9cc;
mem_array[7200] = 16'h3eed;
mem_array[7203] = 16'hec97;
mem_array[7202] = 16'h3e81;
mem_array[7205] = 16'hb650;
mem_array[7204] = 16'h3ee5;
mem_array[7207] = 16'hc0ff;
mem_array[7206] = 16'hbe32;
mem_array[7209] = 16'h26af;
mem_array[7208] = 16'h3f71;
mem_array[7211] = 16'h07cf;
mem_array[7210] = 16'hbf61;
mem_array[7213] = 16'h4a0f;
mem_array[7212] = 16'h3f69;
mem_array[7215] = 16'h9145;
mem_array[7214] = 16'h3d70;
mem_array[7217] = 16'h9151;
mem_array[7216] = 16'h3f23;
mem_array[7219] = 16'h9214;
mem_array[7218] = 16'hbe26;
mem_array[7221] = 16'hf83c;
mem_array[7220] = 16'hbd86;
mem_array[7223] = 16'h5781;
mem_array[7222] = 16'h3aa6;
mem_array[7225] = 16'hdaaf;
mem_array[7224] = 16'h3ea8;
mem_array[7227] = 16'h9a99;
mem_array[7226] = 16'h3dd5;
mem_array[7229] = 16'h76e1;
mem_array[7228] = 16'hbeee;
mem_array[7231] = 16'h50fd;
mem_array[7230] = 16'h3ea4;
mem_array[7233] = 16'hd651;
mem_array[7232] = 16'h3e45;
mem_array[7235] = 16'h2d70;
mem_array[7234] = 16'hbe8a;
mem_array[7237] = 16'h50b2;
mem_array[7236] = 16'hbeea;
mem_array[7239] = 16'h3fa9;
mem_array[7238] = 16'h3d90;
mem_array[7241] = 16'hf054;
mem_array[7240] = 16'hbe65;
mem_array[7243] = 16'he60f;
mem_array[7242] = 16'h3ea5;
mem_array[7245] = 16'h721f;
mem_array[7244] = 16'hbeb1;
mem_array[7247] = 16'h3d75;
mem_array[7246] = 16'h3ed7;
mem_array[7249] = 16'heaf5;
mem_array[7248] = 16'h3eb1;
mem_array[7251] = 16'h0d6b;
mem_array[7250] = 16'hbe2f;
mem_array[7253] = 16'h1772;
mem_array[7252] = 16'h3d83;
mem_array[7255] = 16'h46f0;
mem_array[7254] = 16'h3eb4;
mem_array[7257] = 16'h7b88;
mem_array[7256] = 16'h3e61;
mem_array[7259] = 16'he51e;
mem_array[7258] = 16'hbf12;
mem_array[7261] = 16'h9ce2;
mem_array[7260] = 16'h3eaf;
mem_array[7263] = 16'h9276;
mem_array[7262] = 16'hbdab;
mem_array[7265] = 16'h8f8f;
mem_array[7264] = 16'h3e25;
mem_array[7267] = 16'h2d53;
mem_array[7266] = 16'hbebc;
mem_array[7269] = 16'h9487;
mem_array[7268] = 16'h3e89;
mem_array[7271] = 16'ha35e;
mem_array[7270] = 16'hbc58;
mem_array[7273] = 16'h9fe8;
mem_array[7272] = 16'h3e78;
mem_array[7275] = 16'h0232;
mem_array[7274] = 16'h3e15;
mem_array[7277] = 16'h9f8a;
mem_array[7276] = 16'hbe89;
mem_array[7279] = 16'ha645;
mem_array[7278] = 16'hbf28;
mem_array[7281] = 16'hdf63;
mem_array[7280] = 16'h3d34;
mem_array[7283] = 16'hd010;
mem_array[7282] = 16'h3d2e;
mem_array[7285] = 16'hceda;
mem_array[7284] = 16'h3eb1;
mem_array[7287] = 16'h08b8;
mem_array[7286] = 16'h3ecc;
mem_array[7289] = 16'hbb8f;
mem_array[7288] = 16'hbe24;
mem_array[7291] = 16'h70ee;
mem_array[7290] = 16'h3ec2;
mem_array[7293] = 16'h3c2f;
mem_array[7292] = 16'h3e0f;
mem_array[7295] = 16'he510;
mem_array[7294] = 16'hbe92;
mem_array[7297] = 16'h1c73;
mem_array[7296] = 16'hbf98;
mem_array[7299] = 16'h5a4d;
mem_array[7298] = 16'hbc60;
mem_array[7301] = 16'hf692;
mem_array[7300] = 16'hbeab;
mem_array[7303] = 16'h4201;
mem_array[7302] = 16'h3ebc;
mem_array[7305] = 16'h570f;
mem_array[7304] = 16'h3ca9;
mem_array[7307] = 16'h0878;
mem_array[7306] = 16'h3f02;
mem_array[7309] = 16'h6123;
mem_array[7308] = 16'h3ecc;
mem_array[7311] = 16'h512e;
mem_array[7310] = 16'hbf40;
mem_array[7313] = 16'ha9e5;
mem_array[7312] = 16'h3d5b;
mem_array[7315] = 16'hba3c;
mem_array[7314] = 16'h3e63;
mem_array[7317] = 16'hdeb2;
mem_array[7316] = 16'h3edf;
mem_array[7319] = 16'he961;
mem_array[7318] = 16'hbe01;
mem_array[7321] = 16'h4a0d;
mem_array[7320] = 16'hbefa;
mem_array[7323] = 16'h1085;
mem_array[7322] = 16'hbf09;
mem_array[7325] = 16'hf288;
mem_array[7324] = 16'hbe86;
mem_array[7327] = 16'h99a6;
mem_array[7326] = 16'hbe88;
mem_array[7329] = 16'h50d5;
mem_array[7328] = 16'hbf7a;
mem_array[7331] = 16'h834a;
mem_array[7330] = 16'h3ed2;
mem_array[7333] = 16'h44e0;
mem_array[7332] = 16'h3f00;
mem_array[7335] = 16'h9b1e;
mem_array[7334] = 16'h3ebb;
mem_array[7337] = 16'hdaab;
mem_array[7336] = 16'hbe2d;
mem_array[7339] = 16'h8239;
mem_array[7338] = 16'h3e4a;
mem_array[7341] = 16'habc0;
mem_array[7340] = 16'hbd94;
mem_array[7343] = 16'h972b;
mem_array[7342] = 16'h3d15;
mem_array[7345] = 16'hdf5d;
mem_array[7344] = 16'h3f03;
mem_array[7347] = 16'h8218;
mem_array[7346] = 16'h3ee9;
mem_array[7349] = 16'hf961;
mem_array[7348] = 16'hbe8e;
mem_array[7351] = 16'h0fac;
mem_array[7350] = 16'h3df6;
mem_array[7353] = 16'h755c;
mem_array[7352] = 16'h3d12;
mem_array[7355] = 16'h0080;
mem_array[7354] = 16'hbd98;
mem_array[7357] = 16'h374e;
mem_array[7356] = 16'hbf3a;
mem_array[7359] = 16'h4bc8;
mem_array[7358] = 16'h3de2;
mem_array[7361] = 16'h9ac7;
mem_array[7360] = 16'hbf18;
mem_array[7363] = 16'h3647;
mem_array[7362] = 16'h3dc9;
mem_array[7365] = 16'hdd3d;
mem_array[7364] = 16'hbf0e;
mem_array[7367] = 16'h31c5;
mem_array[7366] = 16'h3d94;
mem_array[7369] = 16'h35c0;
mem_array[7368] = 16'h3e3d;
mem_array[7371] = 16'hc298;
mem_array[7370] = 16'hbf1d;
mem_array[7373] = 16'h1bc2;
mem_array[7372] = 16'h3e88;
mem_array[7375] = 16'h5ebe;
mem_array[7374] = 16'hbe29;
mem_array[7377] = 16'hc7ef;
mem_array[7376] = 16'h3e68;
mem_array[7379] = 16'hfd28;
mem_array[7378] = 16'hbe82;
mem_array[7381] = 16'hc9fc;
mem_array[7380] = 16'hbecd;
mem_array[7383] = 16'hda00;
mem_array[7382] = 16'hbeba;
mem_array[7385] = 16'hec8f;
mem_array[7384] = 16'hbece;
mem_array[7387] = 16'h7904;
mem_array[7386] = 16'h3dee;
mem_array[7389] = 16'h6186;
mem_array[7388] = 16'hbf60;
mem_array[7391] = 16'h398b;
mem_array[7390] = 16'h3ecd;
mem_array[7393] = 16'h95e3;
mem_array[7392] = 16'h3ef6;
mem_array[7395] = 16'heaec;
mem_array[7394] = 16'h3e3b;
mem_array[7397] = 16'hf5e6;
mem_array[7396] = 16'h3eb6;
mem_array[7399] = 16'hbdf0;
mem_array[7398] = 16'h3eb0;
mem_array[7401] = 16'h60b8;
mem_array[7400] = 16'h3b5a;
mem_array[7403] = 16'h3e18;
mem_array[7402] = 16'h3d89;
mem_array[7405] = 16'h7551;
mem_array[7404] = 16'h3ea8;
mem_array[7407] = 16'h8eae;
mem_array[7406] = 16'h3e9d;
mem_array[7409] = 16'hef7c;
mem_array[7408] = 16'hbe7d;
mem_array[7411] = 16'he811;
mem_array[7410] = 16'h3e1c;
mem_array[7413] = 16'h3e78;
mem_array[7412] = 16'h3f0d;
mem_array[7415] = 16'hc9f0;
mem_array[7414] = 16'h3e69;
mem_array[7417] = 16'h95ae;
mem_array[7416] = 16'hbe82;
mem_array[7419] = 16'ha56d;
mem_array[7418] = 16'h3e86;
mem_array[7421] = 16'h5c80;
mem_array[7420] = 16'hbf12;
mem_array[7423] = 16'h2c82;
mem_array[7422] = 16'h3e18;
mem_array[7425] = 16'hac53;
mem_array[7424] = 16'hbf44;
mem_array[7427] = 16'h444e;
mem_array[7426] = 16'hbe13;
mem_array[7429] = 16'h468b;
mem_array[7428] = 16'h3eb9;
mem_array[7431] = 16'hc642;
mem_array[7430] = 16'h3e1c;
mem_array[7433] = 16'h5f4a;
mem_array[7432] = 16'h3eba;
mem_array[7435] = 16'h9143;
mem_array[7434] = 16'hbeaf;
mem_array[7437] = 16'h2a93;
mem_array[7436] = 16'h3ede;
mem_array[7439] = 16'h3c2f;
mem_array[7438] = 16'hbf1c;
mem_array[7441] = 16'hbdfb;
mem_array[7440] = 16'hbea7;
mem_array[7443] = 16'h1c3f;
mem_array[7442] = 16'hbe70;
mem_array[7445] = 16'h2345;
mem_array[7444] = 16'hbda7;
mem_array[7447] = 16'hb6e7;
mem_array[7446] = 16'hbe2f;
mem_array[7449] = 16'hd0a3;
mem_array[7448] = 16'hbf3f;
mem_array[7451] = 16'h0aa3;
mem_array[7450] = 16'hbe15;
mem_array[7453] = 16'h5cf7;
mem_array[7452] = 16'h3edc;
mem_array[7455] = 16'hebcf;
mem_array[7454] = 16'h3e36;
mem_array[7457] = 16'he130;
mem_array[7456] = 16'hbe3d;
mem_array[7459] = 16'hc206;
mem_array[7458] = 16'h3cf8;
mem_array[7461] = 16'h2da8;
mem_array[7460] = 16'h3d3e;
mem_array[7463] = 16'hb1b7;
mem_array[7462] = 16'hbce7;
mem_array[7465] = 16'h387b;
mem_array[7464] = 16'h3c20;
mem_array[7467] = 16'hb09b;
mem_array[7466] = 16'h3f20;
mem_array[7469] = 16'hd355;
mem_array[7468] = 16'hbe58;
mem_array[7471] = 16'ha23e;
mem_array[7470] = 16'h3e94;
mem_array[7473] = 16'haaf8;
mem_array[7472] = 16'h3f07;
mem_array[7475] = 16'hc489;
mem_array[7474] = 16'h3e2d;
mem_array[7477] = 16'h6888;
mem_array[7476] = 16'hbcbd;
mem_array[7479] = 16'h165c;
mem_array[7478] = 16'h3ee2;
mem_array[7481] = 16'h3da0;
mem_array[7480] = 16'hbf09;
mem_array[7483] = 16'heada;
mem_array[7482] = 16'h3e33;
mem_array[7485] = 16'h9bc2;
mem_array[7484] = 16'hbeea;
mem_array[7487] = 16'hcc34;
mem_array[7486] = 16'hbb5a;
mem_array[7489] = 16'hebd3;
mem_array[7488] = 16'h3ce4;
mem_array[7491] = 16'h8eb8;
mem_array[7490] = 16'hbe41;
mem_array[7493] = 16'h8823;
mem_array[7492] = 16'h3e6f;
mem_array[7495] = 16'hcbc9;
mem_array[7494] = 16'hbeff;
mem_array[7497] = 16'h6a86;
mem_array[7496] = 16'h3e1a;
mem_array[7499] = 16'h5cfe;
mem_array[7498] = 16'hbf0c;
mem_array[7501] = 16'hb7e9;
mem_array[7500] = 16'hbf79;
mem_array[7503] = 16'ha880;
mem_array[7502] = 16'hbe5b;
mem_array[7505] = 16'h2aa3;
mem_array[7504] = 16'h3ec7;
mem_array[7507] = 16'h3f92;
mem_array[7506] = 16'h3e14;
mem_array[7509] = 16'h87df;
mem_array[7508] = 16'hbe8c;
mem_array[7511] = 16'h28c4;
mem_array[7510] = 16'hbe06;
mem_array[7513] = 16'h4690;
mem_array[7512] = 16'h3e21;
mem_array[7515] = 16'hb9f9;
mem_array[7514] = 16'h3e49;
mem_array[7517] = 16'hb1f0;
mem_array[7516] = 16'hbf78;
mem_array[7519] = 16'h0492;
mem_array[7518] = 16'h3de6;
mem_array[7521] = 16'hfc00;
mem_array[7520] = 16'hbca8;
mem_array[7523] = 16'h1d51;
mem_array[7522] = 16'hbd11;
mem_array[7525] = 16'h9406;
mem_array[7524] = 16'h3d93;
mem_array[7527] = 16'ha9e6;
mem_array[7526] = 16'h3e42;
mem_array[7529] = 16'h844a;
mem_array[7528] = 16'hbe99;
mem_array[7531] = 16'h5c2f;
mem_array[7530] = 16'h3e68;
mem_array[7533] = 16'h32d2;
mem_array[7532] = 16'hbd21;
mem_array[7535] = 16'h6cd2;
mem_array[7534] = 16'h3e21;
mem_array[7537] = 16'h5d15;
mem_array[7536] = 16'hbf14;
mem_array[7539] = 16'h0d7d;
mem_array[7538] = 16'hbd47;
mem_array[7541] = 16'hf62b;
mem_array[7540] = 16'h3d2f;
mem_array[7543] = 16'hd1b1;
mem_array[7542] = 16'hbd3c;
mem_array[7545] = 16'hbd24;
mem_array[7544] = 16'hbefc;
mem_array[7547] = 16'h2051;
mem_array[7546] = 16'hbdd1;
mem_array[7549] = 16'h5c89;
mem_array[7548] = 16'hbe9c;
mem_array[7551] = 16'h661e;
mem_array[7550] = 16'hbeec;
mem_array[7553] = 16'h6677;
mem_array[7552] = 16'h3df4;
mem_array[7555] = 16'h8fe6;
mem_array[7554] = 16'hbe4a;
mem_array[7557] = 16'hd9b6;
mem_array[7556] = 16'h3deb;
mem_array[7559] = 16'h542c;
mem_array[7558] = 16'hbebc;
mem_array[7561] = 16'he7fd;
mem_array[7560] = 16'h3d5e;
mem_array[7563] = 16'hacf8;
mem_array[7562] = 16'hbea5;
mem_array[7565] = 16'h4a4e;
mem_array[7564] = 16'h3e32;
mem_array[7567] = 16'hd7c1;
mem_array[7566] = 16'h3b92;
mem_array[7569] = 16'ha2e5;
mem_array[7568] = 16'h3d35;
mem_array[7571] = 16'h3e50;
mem_array[7570] = 16'h3d83;
mem_array[7573] = 16'h485f;
mem_array[7572] = 16'hbc0e;
mem_array[7575] = 16'h349d;
mem_array[7574] = 16'h3e41;
mem_array[7577] = 16'heffb;
mem_array[7576] = 16'hbf7a;
mem_array[7579] = 16'hab35;
mem_array[7578] = 16'h3c3b;
mem_array[7581] = 16'h7f70;
mem_array[7580] = 16'h3d5b;
mem_array[7583] = 16'hf7f4;
mem_array[7582] = 16'h3db9;
mem_array[7585] = 16'hc341;
mem_array[7584] = 16'h3e43;
mem_array[7587] = 16'hac9b;
mem_array[7586] = 16'h3e38;
mem_array[7589] = 16'h768e;
mem_array[7588] = 16'hbdf0;
mem_array[7591] = 16'hbee9;
mem_array[7590] = 16'h3e19;
mem_array[7593] = 16'h4d3c;
mem_array[7592] = 16'h3dac;
mem_array[7595] = 16'h7149;
mem_array[7594] = 16'hbf35;
mem_array[7597] = 16'hd8e0;
mem_array[7596] = 16'hbfb8;
mem_array[7599] = 16'h9140;
mem_array[7598] = 16'h3e9e;
mem_array[7601] = 16'hc9d2;
mem_array[7600] = 16'hbb62;
mem_array[7603] = 16'h4605;
mem_array[7602] = 16'h3da6;
mem_array[7605] = 16'h289b;
mem_array[7604] = 16'hbe87;
mem_array[7607] = 16'h940b;
mem_array[7606] = 16'hbe0b;
mem_array[7609] = 16'h4936;
mem_array[7608] = 16'hbe48;
mem_array[7611] = 16'h703a;
mem_array[7610] = 16'h3ee8;
mem_array[7613] = 16'h1f87;
mem_array[7612] = 16'h3e9a;
mem_array[7615] = 16'ha1f5;
mem_array[7614] = 16'hbe53;
mem_array[7617] = 16'haaa3;
mem_array[7616] = 16'h3e6a;
mem_array[7619] = 16'h9381;
mem_array[7618] = 16'hbed6;
mem_array[7621] = 16'h653a;
mem_array[7620] = 16'h3f5d;
mem_array[7623] = 16'h04f3;
mem_array[7622] = 16'hbf10;
mem_array[7625] = 16'hb8f5;
mem_array[7624] = 16'hbd00;
mem_array[7627] = 16'h152e;
mem_array[7626] = 16'h3d04;
mem_array[7629] = 16'h9a5b;
mem_array[7628] = 16'hbefd;
mem_array[7631] = 16'h5dea;
mem_array[7630] = 16'h3dd5;
mem_array[7633] = 16'hb2bb;
mem_array[7632] = 16'h3da7;
mem_array[7635] = 16'h7450;
mem_array[7634] = 16'h3e49;
mem_array[7637] = 16'hf8ac;
mem_array[7636] = 16'hbf22;
mem_array[7639] = 16'h4c6b;
mem_array[7638] = 16'h3e11;
mem_array[7641] = 16'h44ce;
mem_array[7640] = 16'hbe1b;
mem_array[7643] = 16'hf6e1;
mem_array[7642] = 16'h3c85;
mem_array[7645] = 16'he79c;
mem_array[7644] = 16'hbde6;
mem_array[7647] = 16'h1905;
mem_array[7646] = 16'h3b86;
mem_array[7649] = 16'h9c38;
mem_array[7648] = 16'h3ded;
mem_array[7651] = 16'haef2;
mem_array[7650] = 16'h3e06;
mem_array[7653] = 16'h2dc4;
mem_array[7652] = 16'hbea2;
mem_array[7655] = 16'h38b8;
mem_array[7654] = 16'hbf7e;
mem_array[7657] = 16'hb9e4;
mem_array[7656] = 16'hbf8c;
mem_array[7659] = 16'hebe2;
mem_array[7658] = 16'hbeb2;
mem_array[7661] = 16'hea35;
mem_array[7660] = 16'hbf1c;
mem_array[7663] = 16'heb74;
mem_array[7662] = 16'h3e4d;
mem_array[7665] = 16'h9f1b;
mem_array[7664] = 16'hbe08;
mem_array[7667] = 16'h21fd;
mem_array[7666] = 16'hbe33;
mem_array[7669] = 16'hc249;
mem_array[7668] = 16'h3d92;
mem_array[7671] = 16'h5f14;
mem_array[7670] = 16'hbe35;
mem_array[7673] = 16'h5fc4;
mem_array[7672] = 16'h3e2d;
mem_array[7675] = 16'h0e2b;
mem_array[7674] = 16'hbe79;
mem_array[7677] = 16'hdcb9;
mem_array[7676] = 16'h3e9a;
mem_array[7679] = 16'ha975;
mem_array[7678] = 16'hbe36;
mem_array[7681] = 16'hd360;
mem_array[7680] = 16'h3e88;
mem_array[7683] = 16'h3a33;
mem_array[7682] = 16'hbd07;
mem_array[7685] = 16'h98ae;
mem_array[7684] = 16'hbe48;
mem_array[7687] = 16'h0468;
mem_array[7686] = 16'h3e6e;
mem_array[7689] = 16'hc0f6;
mem_array[7688] = 16'hbf3c;
mem_array[7691] = 16'he3bc;
mem_array[7690] = 16'h3c0c;
mem_array[7693] = 16'h5cb7;
mem_array[7692] = 16'h3e10;
mem_array[7695] = 16'hf71a;
mem_array[7694] = 16'hbc1a;
mem_array[7697] = 16'h238d;
mem_array[7696] = 16'h3d8c;
mem_array[7699] = 16'hec4e;
mem_array[7698] = 16'hbe23;
mem_array[7701] = 16'h7069;
mem_array[7700] = 16'h3c9c;
mem_array[7703] = 16'hbf3b;
mem_array[7702] = 16'hbd8e;
mem_array[7705] = 16'h473e;
mem_array[7704] = 16'hbea9;
mem_array[7707] = 16'h42d3;
mem_array[7706] = 16'hbd65;
mem_array[7709] = 16'h0385;
mem_array[7708] = 16'h3e05;
mem_array[7711] = 16'h0acb;
mem_array[7710] = 16'h3e21;
mem_array[7713] = 16'haaf9;
mem_array[7712] = 16'h3e90;
mem_array[7715] = 16'h28bf;
mem_array[7714] = 16'h3cf9;
mem_array[7717] = 16'hef33;
mem_array[7716] = 16'h3c29;
mem_array[7719] = 16'hd1c2;
mem_array[7718] = 16'hbeca;
mem_array[7721] = 16'hf2de;
mem_array[7720] = 16'hbceb;
mem_array[7723] = 16'h9d4c;
mem_array[7722] = 16'h3e7a;
mem_array[7725] = 16'hcc36;
mem_array[7724] = 16'hbe20;
mem_array[7727] = 16'hbbbf;
mem_array[7726] = 16'hbdd0;
mem_array[7729] = 16'h4436;
mem_array[7728] = 16'hbe00;
mem_array[7731] = 16'h9777;
mem_array[7730] = 16'hbeaf;
mem_array[7733] = 16'h0910;
mem_array[7732] = 16'h3d9e;
mem_array[7735] = 16'h879d;
mem_array[7734] = 16'hbdd9;
mem_array[7737] = 16'hb6e3;
mem_array[7736] = 16'h3edb;
mem_array[7739] = 16'hedca;
mem_array[7738] = 16'h3e38;
mem_array[7741] = 16'he441;
mem_array[7740] = 16'h3e1f;
mem_array[7743] = 16'h9832;
mem_array[7742] = 16'hbe4c;
mem_array[7745] = 16'h2b02;
mem_array[7744] = 16'hbe7f;
mem_array[7747] = 16'hac25;
mem_array[7746] = 16'hbd8e;
mem_array[7749] = 16'h8479;
mem_array[7748] = 16'hbf4f;
mem_array[7751] = 16'h8878;
mem_array[7750] = 16'hbd62;
mem_array[7753] = 16'h2771;
mem_array[7752] = 16'h3e24;
mem_array[7755] = 16'h9b5d;
mem_array[7754] = 16'hbe84;
mem_array[7757] = 16'h9196;
mem_array[7756] = 16'h3e8f;
mem_array[7759] = 16'he7f0;
mem_array[7758] = 16'h3e52;
mem_array[7761] = 16'h46ea;
mem_array[7760] = 16'hbda4;
mem_array[7763] = 16'he170;
mem_array[7762] = 16'h3bd2;
mem_array[7765] = 16'hb298;
mem_array[7764] = 16'hbe74;
mem_array[7767] = 16'h0441;
mem_array[7766] = 16'h3e87;
mem_array[7769] = 16'h7604;
mem_array[7768] = 16'hbe0c;
mem_array[7771] = 16'h9a92;
mem_array[7770] = 16'h3dc5;
mem_array[7773] = 16'h09ea;
mem_array[7772] = 16'hbd00;
mem_array[7775] = 16'he1e3;
mem_array[7774] = 16'hbefa;
mem_array[7777] = 16'h4b28;
mem_array[7776] = 16'hbeeb;
mem_array[7779] = 16'h7cd5;
mem_array[7778] = 16'hbda9;
mem_array[7781] = 16'h889e;
mem_array[7780] = 16'h3cbf;
mem_array[7783] = 16'hd4b4;
mem_array[7782] = 16'h3e89;
mem_array[7785] = 16'hbb41;
mem_array[7784] = 16'h3e4d;
mem_array[7787] = 16'h47d5;
mem_array[7786] = 16'h3e0f;
mem_array[7789] = 16'h9b64;
mem_array[7788] = 16'h3d27;
mem_array[7791] = 16'heb42;
mem_array[7790] = 16'h3d80;
mem_array[7793] = 16'h7f42;
mem_array[7792] = 16'h3e12;
mem_array[7795] = 16'hc8f1;
mem_array[7794] = 16'h3e2f;
mem_array[7797] = 16'hd80e;
mem_array[7796] = 16'h3f08;
mem_array[7799] = 16'h48df;
mem_array[7798] = 16'hbe86;
mem_array[7801] = 16'he81b;
mem_array[7800] = 16'h3e5a;
mem_array[7803] = 16'h8b01;
mem_array[7802] = 16'hbeb3;
mem_array[7805] = 16'h207e;
mem_array[7804] = 16'hbdfa;
mem_array[7807] = 16'ha15f;
mem_array[7806] = 16'h3eeb;
mem_array[7809] = 16'hb0b9;
mem_array[7808] = 16'hbe75;
mem_array[7811] = 16'h436f;
mem_array[7810] = 16'h3ec8;
mem_array[7813] = 16'h701d;
mem_array[7812] = 16'h3dd1;
mem_array[7815] = 16'hc901;
mem_array[7814] = 16'hbd61;
mem_array[7817] = 16'ha92b;
mem_array[7816] = 16'hbdba;
mem_array[7819] = 16'h4173;
mem_array[7818] = 16'h3dd8;
mem_array[7821] = 16'h9524;
mem_array[7820] = 16'hbcc4;
mem_array[7823] = 16'hd8b5;
mem_array[7822] = 16'hbdd0;
mem_array[7825] = 16'hb93c;
mem_array[7824] = 16'h3c54;
mem_array[7827] = 16'hdb20;
mem_array[7826] = 16'h3e94;
mem_array[7829] = 16'h6fd4;
mem_array[7828] = 16'h3d87;
mem_array[7831] = 16'hf8cd;
mem_array[7830] = 16'hbe9a;
mem_array[7833] = 16'h20f3;
mem_array[7832] = 16'hbe0c;
mem_array[7835] = 16'h0ff8;
mem_array[7834] = 16'hbe66;
mem_array[7837] = 16'h6071;
mem_array[7836] = 16'hbebc;
mem_array[7839] = 16'h59ae;
mem_array[7838] = 16'hbef9;
mem_array[7841] = 16'h7778;
mem_array[7840] = 16'hbecc;
mem_array[7843] = 16'h782a;
mem_array[7842] = 16'hbb56;
mem_array[7845] = 16'h81f8;
mem_array[7844] = 16'hbed8;
mem_array[7847] = 16'h3ad0;
mem_array[7846] = 16'hbd41;
mem_array[7849] = 16'h62e0;
mem_array[7848] = 16'h3d91;
mem_array[7851] = 16'h56fc;
mem_array[7850] = 16'hbf83;
mem_array[7853] = 16'hce35;
mem_array[7852] = 16'h3b7b;
mem_array[7855] = 16'h2737;
mem_array[7854] = 16'hbde7;
mem_array[7857] = 16'h59d7;
mem_array[7856] = 16'h3e95;
mem_array[7859] = 16'h2182;
mem_array[7858] = 16'hbbfc;
mem_array[7861] = 16'hf4a3;
mem_array[7860] = 16'h3f0c;
mem_array[7863] = 16'ha1c3;
mem_array[7862] = 16'h3eb3;
mem_array[7865] = 16'h6c3c;
mem_array[7864] = 16'hbea3;
mem_array[7867] = 16'he93f;
mem_array[7866] = 16'h3d70;
mem_array[7869] = 16'hd9ad;
mem_array[7868] = 16'h3eb7;
mem_array[7871] = 16'h4451;
mem_array[7870] = 16'h3d29;
mem_array[7873] = 16'h73c5;
mem_array[7872] = 16'hbe3c;
mem_array[7875] = 16'h6fde;
mem_array[7874] = 16'hbe28;
mem_array[7877] = 16'h492e;
mem_array[7876] = 16'hbe30;
mem_array[7879] = 16'h7bad;
mem_array[7878] = 16'hbf02;
mem_array[7881] = 16'h8101;
mem_array[7880] = 16'hbc13;
mem_array[7883] = 16'h1642;
mem_array[7882] = 16'h3c94;
mem_array[7885] = 16'hc67d;
mem_array[7884] = 16'hbed3;
mem_array[7887] = 16'h1d9e;
mem_array[7886] = 16'h3e36;
mem_array[7889] = 16'hb77a;
mem_array[7888] = 16'hbdee;
mem_array[7891] = 16'ha858;
mem_array[7890] = 16'h3cc1;
mem_array[7893] = 16'hb92a;
mem_array[7892] = 16'h3ee2;
mem_array[7895] = 16'h89e7;
mem_array[7894] = 16'hbdba;
mem_array[7897] = 16'h59cb;
mem_array[7896] = 16'h3eef;
mem_array[7899] = 16'hf6e2;
mem_array[7898] = 16'hbd48;
mem_array[7901] = 16'hc29d;
mem_array[7900] = 16'h3ed9;
mem_array[7903] = 16'h54f4;
mem_array[7902] = 16'hbe93;
mem_array[7905] = 16'hca3e;
mem_array[7904] = 16'h3e50;
mem_array[7907] = 16'h25a6;
mem_array[7906] = 16'hbe7f;
mem_array[7909] = 16'h2a61;
mem_array[7908] = 16'hbd99;
mem_array[7911] = 16'h56ca;
mem_array[7910] = 16'hbe52;
mem_array[7913] = 16'hb7f6;
mem_array[7912] = 16'h3cf4;
mem_array[7915] = 16'h8bc3;
mem_array[7914] = 16'hbe8d;
mem_array[7917] = 16'h5f84;
mem_array[7916] = 16'h3d5e;
mem_array[7919] = 16'hd1eb;
mem_array[7918] = 16'h3d92;
mem_array[7921] = 16'hc96c;
mem_array[7920] = 16'h3f33;
mem_array[7923] = 16'hffd8;
mem_array[7922] = 16'h3d31;
mem_array[7925] = 16'hc863;
mem_array[7924] = 16'h3e90;
mem_array[7927] = 16'h701c;
mem_array[7926] = 16'hbe4d;
mem_array[7929] = 16'haac1;
mem_array[7928] = 16'h3f2a;
mem_array[7931] = 16'h06f9;
mem_array[7930] = 16'hbe6e;
mem_array[7933] = 16'he92b;
mem_array[7932] = 16'hbec4;
mem_array[7935] = 16'h18da;
mem_array[7934] = 16'hbc98;
mem_array[7937] = 16'h1f62;
mem_array[7936] = 16'hbe98;
mem_array[7939] = 16'h14ec;
mem_array[7938] = 16'hbf40;
mem_array[7941] = 16'h2a68;
mem_array[7940] = 16'h3dac;
mem_array[7943] = 16'h57dc;
mem_array[7942] = 16'hbcce;
mem_array[7945] = 16'h6570;
mem_array[7944] = 16'hbed9;
mem_array[7947] = 16'hb012;
mem_array[7946] = 16'hbd78;
mem_array[7949] = 16'h0a3a;
mem_array[7948] = 16'h3dcc;
mem_array[7951] = 16'h7683;
mem_array[7950] = 16'h3e0e;
mem_array[7953] = 16'h0a0e;
mem_array[7952] = 16'h3de1;
mem_array[7955] = 16'h2059;
mem_array[7954] = 16'hbda3;
mem_array[7957] = 16'hf6c0;
mem_array[7956] = 16'h3e8d;
mem_array[7959] = 16'h5e88;
mem_array[7958] = 16'h3e63;
mem_array[7961] = 16'h2ac9;
mem_array[7960] = 16'h3e2f;
mem_array[7963] = 16'h26f5;
mem_array[7962] = 16'hbc1c;
mem_array[7965] = 16'h888b;
mem_array[7964] = 16'h3edf;
mem_array[7967] = 16'hb8b3;
mem_array[7966] = 16'hbd3e;
mem_array[7969] = 16'h2ba4;
mem_array[7968] = 16'h3d0b;
mem_array[7971] = 16'h5988;
mem_array[7970] = 16'hbedb;
mem_array[7973] = 16'h54ab;
mem_array[7972] = 16'h3e26;
mem_array[7975] = 16'hc737;
mem_array[7974] = 16'hbe14;
mem_array[7977] = 16'hf1e1;
mem_array[7976] = 16'h3d08;
mem_array[7979] = 16'h5cf0;
mem_array[7978] = 16'h3e1e;
mem_array[7981] = 16'had68;
mem_array[7980] = 16'hbdc9;
mem_array[7983] = 16'hff85;
mem_array[7982] = 16'h3dee;
mem_array[7985] = 16'h1e4b;
mem_array[7984] = 16'hbe44;
mem_array[7987] = 16'h5411;
mem_array[7986] = 16'h3d9a;
mem_array[7989] = 16'h3b4d;
mem_array[7988] = 16'h3f86;
mem_array[7991] = 16'hee2b;
mem_array[7990] = 16'h3e5f;
mem_array[7993] = 16'h4428;
mem_array[7992] = 16'hbf01;
mem_array[7995] = 16'h9538;
mem_array[7994] = 16'h3d3e;
mem_array[7997] = 16'h4ac0;
mem_array[7996] = 16'hbee7;
mem_array[7999] = 16'h6707;
mem_array[7998] = 16'hbf29;
mem_array[8001] = 16'hb34b;
mem_array[8000] = 16'hbd96;
mem_array[8003] = 16'hf16e;
mem_array[8002] = 16'hbd1c;
mem_array[8005] = 16'h1d28;
mem_array[8004] = 16'hbb89;
mem_array[8007] = 16'heb58;
mem_array[8006] = 16'hbeab;
mem_array[8009] = 16'hbd41;
mem_array[8008] = 16'hbe49;
mem_array[8011] = 16'h3e56;
mem_array[8010] = 16'h3c3e;
mem_array[8013] = 16'h3750;
mem_array[8012] = 16'hbf29;
mem_array[8015] = 16'hfad4;
mem_array[8014] = 16'h3f19;
mem_array[8017] = 16'h721d;
mem_array[8016] = 16'h3e75;
mem_array[8019] = 16'h8413;
mem_array[8018] = 16'h3ec7;
mem_array[8021] = 16'h998f;
mem_array[8020] = 16'h3ea3;
mem_array[8023] = 16'h0b3f;
mem_array[8022] = 16'h3f08;
mem_array[8025] = 16'hd3e0;
mem_array[8024] = 16'hbded;
mem_array[8027] = 16'hed84;
mem_array[8026] = 16'h3e28;
mem_array[8029] = 16'hf980;
mem_array[8028] = 16'hbece;
mem_array[8031] = 16'hed8a;
mem_array[8030] = 16'hbebc;
mem_array[8033] = 16'h949c;
mem_array[8032] = 16'h3ec7;
mem_array[8035] = 16'h372a;
mem_array[8034] = 16'h3da8;
mem_array[8037] = 16'h468a;
mem_array[8036] = 16'hbd27;
mem_array[8039] = 16'h6806;
mem_array[8038] = 16'h3ef3;
mem_array[8041] = 16'h921d;
mem_array[8040] = 16'h3ee4;
mem_array[8043] = 16'hfec1;
mem_array[8042] = 16'hbe2f;
mem_array[8045] = 16'h43ea;
mem_array[8044] = 16'hbe25;
mem_array[8047] = 16'h53f5;
mem_array[8046] = 16'h3e1b;
mem_array[8049] = 16'h3959;
mem_array[8048] = 16'h3f9e;
mem_array[8051] = 16'hd538;
mem_array[8050] = 16'h3ec2;
mem_array[8053] = 16'h388b;
mem_array[8052] = 16'hbece;
mem_array[8055] = 16'h45aa;
mem_array[8054] = 16'hbdcc;
mem_array[8057] = 16'h4574;
mem_array[8056] = 16'hbefe;
mem_array[8059] = 16'h2cf9;
mem_array[8058] = 16'hbebf;
mem_array[8061] = 16'hecb0;
mem_array[8060] = 16'hbd15;
mem_array[8063] = 16'hc572;
mem_array[8062] = 16'h3cac;
mem_array[8065] = 16'h1582;
mem_array[8064] = 16'hbd77;
mem_array[8067] = 16'h76ec;
mem_array[8066] = 16'h3eab;
mem_array[8069] = 16'h90d4;
mem_array[8068] = 16'h3e8c;
mem_array[8071] = 16'h261d;
mem_array[8070] = 16'hbe3f;
mem_array[8073] = 16'h11f7;
mem_array[8072] = 16'hbe2f;
mem_array[8075] = 16'hde3d;
mem_array[8074] = 16'h3f60;
mem_array[8077] = 16'h7b42;
mem_array[8076] = 16'hbc70;
mem_array[8079] = 16'hdc3c;
mem_array[8078] = 16'h3f52;
mem_array[8081] = 16'hf335;
mem_array[8080] = 16'hbed1;
mem_array[8083] = 16'h3f0c;
mem_array[8082] = 16'h3db3;
mem_array[8085] = 16'h7ade;
mem_array[8084] = 16'h3de9;
mem_array[8087] = 16'h7250;
mem_array[8086] = 16'h3e5a;
mem_array[8089] = 16'h9f39;
mem_array[8088] = 16'h3f03;
mem_array[8091] = 16'h1a79;
mem_array[8090] = 16'hbeed;
mem_array[8093] = 16'h94a0;
mem_array[8092] = 16'h3efa;
mem_array[8095] = 16'hfa00;
mem_array[8094] = 16'h3e19;
mem_array[8097] = 16'h4c22;
mem_array[8096] = 16'hbeba;
mem_array[8099] = 16'hb8cc;
mem_array[8098] = 16'h3e78;
mem_array[8101] = 16'h1c2c;
mem_array[8100] = 16'h3cb8;
mem_array[8103] = 16'ha404;
mem_array[8102] = 16'h3e35;
mem_array[8105] = 16'h1d88;
mem_array[8104] = 16'h3f16;
mem_array[8107] = 16'h6f07;
mem_array[8106] = 16'hbe2d;
mem_array[8109] = 16'h9f2d;
mem_array[8108] = 16'h3f5c;
mem_array[8111] = 16'h579a;
mem_array[8110] = 16'h3f0f;
mem_array[8113] = 16'hafd2;
mem_array[8112] = 16'hbec2;
mem_array[8115] = 16'he17a;
mem_array[8114] = 16'hbe83;
mem_array[8117] = 16'h390e;
mem_array[8116] = 16'hbed8;
mem_array[8119] = 16'hd9e6;
mem_array[8118] = 16'hbf12;
mem_array[8121] = 16'he5d1;
mem_array[8120] = 16'h3b34;
mem_array[8123] = 16'h6256;
mem_array[8122] = 16'h3ccf;
mem_array[8125] = 16'hb939;
mem_array[8124] = 16'h3d88;
mem_array[8127] = 16'h6714;
mem_array[8126] = 16'hbf34;
mem_array[8129] = 16'hcca3;
mem_array[8128] = 16'hbf0a;
mem_array[8131] = 16'h0ad6;
mem_array[8130] = 16'hbe71;
mem_array[8133] = 16'h3102;
mem_array[8132] = 16'hbea4;
mem_array[8135] = 16'hd751;
mem_array[8134] = 16'hbe4a;
mem_array[8137] = 16'hf6bd;
mem_array[8136] = 16'h3e7f;
mem_array[8139] = 16'h43de;
mem_array[8138] = 16'h3f24;
mem_array[8141] = 16'h6082;
mem_array[8140] = 16'h3f26;
mem_array[8143] = 16'ha9a3;
mem_array[8142] = 16'h3ec1;
mem_array[8145] = 16'h35cd;
mem_array[8144] = 16'hbe06;
mem_array[8147] = 16'h4258;
mem_array[8146] = 16'h3eb2;
mem_array[8149] = 16'hdcae;
mem_array[8148] = 16'hbf6c;
mem_array[8151] = 16'h4090;
mem_array[8150] = 16'h3d87;
mem_array[8153] = 16'h09d5;
mem_array[8152] = 16'h3f21;
mem_array[8155] = 16'h33ce;
mem_array[8154] = 16'h3eb9;
mem_array[8157] = 16'h7027;
mem_array[8156] = 16'hbe86;
mem_array[8159] = 16'ha87b;
mem_array[8158] = 16'h3e12;
mem_array[8161] = 16'hd23c;
mem_array[8160] = 16'hbf15;
mem_array[8163] = 16'h0751;
mem_array[8162] = 16'h3ee1;
mem_array[8165] = 16'hc4c7;
mem_array[8164] = 16'hbeb9;
mem_array[8167] = 16'hf70c;
mem_array[8166] = 16'hbe53;
mem_array[8169] = 16'h175f;
mem_array[8168] = 16'hbd11;
mem_array[8171] = 16'h74c1;
mem_array[8170] = 16'h3ea2;
mem_array[8173] = 16'h933f;
mem_array[8172] = 16'hbeaa;
mem_array[8175] = 16'h341a;
mem_array[8174] = 16'hbd57;
mem_array[8177] = 16'hf0f6;
mem_array[8176] = 16'hbed1;
mem_array[8179] = 16'h96b6;
mem_array[8178] = 16'hbe35;
mem_array[8181] = 16'h0cb8;
mem_array[8180] = 16'hbd0a;
mem_array[8183] = 16'hb9b0;
mem_array[8182] = 16'h3c22;
mem_array[8185] = 16'h3205;
mem_array[8184] = 16'hbe37;
mem_array[8187] = 16'hd716;
mem_array[8186] = 16'hbfab;
mem_array[8189] = 16'ha1a9;
mem_array[8188] = 16'hbfbd;
mem_array[8191] = 16'hac9b;
mem_array[8190] = 16'hbf31;
mem_array[8193] = 16'h8f48;
mem_array[8192] = 16'hbf2a;
mem_array[8195] = 16'h40ad;
mem_array[8194] = 16'hbe8c;
mem_array[8197] = 16'hb3e9;
mem_array[8196] = 16'hbe99;
mem_array[8199] = 16'hd15e;
mem_array[8198] = 16'h3ead;
mem_array[8201] = 16'hacbb;
mem_array[8200] = 16'h3ed5;
mem_array[8203] = 16'h3899;
mem_array[8202] = 16'h3f75;
mem_array[8205] = 16'h8f19;
mem_array[8204] = 16'hbfc1;
mem_array[8207] = 16'h7324;
mem_array[8206] = 16'h3eab;
mem_array[8209] = 16'hfa30;
mem_array[8208] = 16'hbedf;
mem_array[8211] = 16'hcf76;
mem_array[8210] = 16'hbd46;
mem_array[8213] = 16'h85f6;
mem_array[8212] = 16'h3f72;
mem_array[8215] = 16'h7030;
mem_array[8214] = 16'h3ee2;
mem_array[8217] = 16'h3a35;
mem_array[8216] = 16'hbefe;
mem_array[8219] = 16'h1a77;
mem_array[8218] = 16'hbe9f;
mem_array[8221] = 16'hb36d;
mem_array[8220] = 16'hbf65;
mem_array[8223] = 16'h3025;
mem_array[8222] = 16'h3f08;
mem_array[8225] = 16'h9fad;
mem_array[8224] = 16'hbf46;
mem_array[8227] = 16'h371f;
mem_array[8226] = 16'hbf04;
mem_array[8229] = 16'h5311;
mem_array[8228] = 16'h3f90;
mem_array[8231] = 16'h2d1a;
mem_array[8230] = 16'h3ed6;
mem_array[8233] = 16'h1975;
mem_array[8232] = 16'h3eea;
mem_array[8235] = 16'he44f;
mem_array[8234] = 16'hbebb;
mem_array[8237] = 16'h15f0;
mem_array[8236] = 16'h3f45;
mem_array[8239] = 16'hfdde;
mem_array[8238] = 16'hbbdc;
mem_array[8241] = 16'hde19;
mem_array[8240] = 16'hbcb1;
mem_array[8243] = 16'hfeca;
mem_array[8242] = 16'hbdd5;
mem_array[8245] = 16'h4e98;
mem_array[8244] = 16'h3e39;
mem_array[8247] = 16'hf71b;
mem_array[8246] = 16'h3e52;
mem_array[8249] = 16'he3b7;
mem_array[8248] = 16'hbf81;
mem_array[8251] = 16'h4fa5;
mem_array[8250] = 16'hbed4;
mem_array[8253] = 16'ha0c9;
mem_array[8252] = 16'hbf93;
mem_array[8255] = 16'hffe1;
mem_array[8254] = 16'h3f09;
mem_array[8257] = 16'h2004;
mem_array[8256] = 16'h3f81;
mem_array[8259] = 16'h284b;
mem_array[8258] = 16'h3f8d;
mem_array[8261] = 16'h0808;
mem_array[8260] = 16'h3e3e;
mem_array[8263] = 16'h9bb7;
mem_array[8262] = 16'h3ef4;
mem_array[8265] = 16'h1f88;
mem_array[8264] = 16'hbed9;
mem_array[8267] = 16'hc532;
mem_array[8266] = 16'hbed3;
mem_array[8269] = 16'h7f02;
mem_array[8268] = 16'hbd41;
mem_array[8271] = 16'h5e8a;
mem_array[8270] = 16'hbd56;
mem_array[8273] = 16'hed5b;
mem_array[8272] = 16'h3f2c;
mem_array[8275] = 16'hdf26;
mem_array[8274] = 16'h3f0c;
mem_array[8277] = 16'h178f;
mem_array[8276] = 16'h3ea4;
mem_array[8279] = 16'h0719;
mem_array[8278] = 16'hbf7a;
mem_array[8281] = 16'h23fd;
mem_array[8280] = 16'hbe75;
mem_array[8283] = 16'h7365;
mem_array[8282] = 16'h3c65;
mem_array[8285] = 16'h33e5;
mem_array[8284] = 16'hbe3f;
mem_array[8287] = 16'hfe78;
mem_array[8286] = 16'hbe9f;
mem_array[8289] = 16'h7bb7;
mem_array[8288] = 16'h3f07;
mem_array[8291] = 16'hba93;
mem_array[8290] = 16'h3f36;
mem_array[8293] = 16'hd617;
mem_array[8292] = 16'hbb36;
mem_array[8295] = 16'h004a;
mem_array[8294] = 16'hbede;
mem_array[8297] = 16'h69ef;
mem_array[8296] = 16'hbcdf;
mem_array[8299] = 16'hdeda;
mem_array[8298] = 16'h3d2d;
mem_array[8301] = 16'h1576;
mem_array[8300] = 16'h3d10;
mem_array[8303] = 16'hb8ce;
mem_array[8302] = 16'hbd2d;
mem_array[8305] = 16'h68be;
mem_array[8304] = 16'h3ea0;
mem_array[8307] = 16'ha2f2;
mem_array[8306] = 16'hbd82;
mem_array[8309] = 16'h9404;
mem_array[8308] = 16'hbe01;
mem_array[8311] = 16'hb00f;
mem_array[8310] = 16'hbcfd;
mem_array[8313] = 16'h7aa6;
mem_array[8312] = 16'hbf05;
mem_array[8315] = 16'hd86f;
mem_array[8314] = 16'h3e50;
mem_array[8317] = 16'h0090;
mem_array[8316] = 16'h3d31;
mem_array[8319] = 16'h9679;
mem_array[8318] = 16'hbc19;
mem_array[8321] = 16'he5c1;
mem_array[8320] = 16'hbe7c;
mem_array[8323] = 16'h16b1;
mem_array[8322] = 16'h3ea3;
mem_array[8325] = 16'hd5fd;
mem_array[8324] = 16'h3d74;
mem_array[8327] = 16'hb702;
mem_array[8326] = 16'hbed6;
mem_array[8329] = 16'hb376;
mem_array[8328] = 16'hbd0d;
mem_array[8331] = 16'h0b1c;
mem_array[8330] = 16'h3c99;
mem_array[8333] = 16'h9161;
mem_array[8332] = 16'h3f4f;
mem_array[8335] = 16'hcdd8;
mem_array[8334] = 16'hbefe;
mem_array[8337] = 16'h7f5e;
mem_array[8336] = 16'hbdd5;
mem_array[8339] = 16'h73ac;
mem_array[8338] = 16'hbf48;
mem_array[8341] = 16'hc625;
mem_array[8340] = 16'hbd4c;
mem_array[8343] = 16'h59f0;
mem_array[8342] = 16'hbda2;
mem_array[8345] = 16'h7c55;
mem_array[8344] = 16'hbe56;
mem_array[8347] = 16'heaa2;
mem_array[8346] = 16'hbd44;
mem_array[8349] = 16'h2710;
mem_array[8348] = 16'hbd8c;
mem_array[8351] = 16'h27ac;
mem_array[8350] = 16'h3e7a;
mem_array[8353] = 16'hf216;
mem_array[8352] = 16'hbcd2;
mem_array[8355] = 16'hd63d;
mem_array[8354] = 16'hbd8e;
mem_array[8357] = 16'h97d7;
mem_array[8356] = 16'h3d99;
mem_array[8359] = 16'h43f1;
mem_array[8358] = 16'hbd7f;
mem_array[8361] = 16'ha9d0;
mem_array[8360] = 16'h3cf9;
mem_array[8363] = 16'h938d;
mem_array[8362] = 16'h3ca2;
mem_array[8365] = 16'h8605;
mem_array[8364] = 16'h3f38;
mem_array[8367] = 16'h889c;
mem_array[8366] = 16'hbe3d;
mem_array[8369] = 16'h1e27;
mem_array[8368] = 16'hbe04;
mem_array[8371] = 16'h1250;
mem_array[8370] = 16'hbebd;
mem_array[8373] = 16'h6eeb;
mem_array[8372] = 16'hbee4;
mem_array[8375] = 16'h73b3;
mem_array[8374] = 16'hbe34;
mem_array[8377] = 16'hf827;
mem_array[8376] = 16'hbd04;
mem_array[8379] = 16'h7562;
mem_array[8378] = 16'hbd8e;
mem_array[8381] = 16'h119f;
mem_array[8380] = 16'hbe91;
mem_array[8383] = 16'h03aa;
mem_array[8382] = 16'hbcb4;
mem_array[8385] = 16'h68ad;
mem_array[8384] = 16'h3d68;
mem_array[8387] = 16'h4838;
mem_array[8386] = 16'h3e9a;
mem_array[8389] = 16'h2071;
mem_array[8388] = 16'hbd56;
mem_array[8391] = 16'h5215;
mem_array[8390] = 16'h3d74;
mem_array[8393] = 16'hb0f3;
mem_array[8392] = 16'hbe23;
mem_array[8395] = 16'hf209;
mem_array[8394] = 16'hbd9a;
mem_array[8397] = 16'h7e63;
mem_array[8396] = 16'hbd0c;
mem_array[8399] = 16'hd4af;
mem_array[8398] = 16'hbdd7;
mem_array[8401] = 16'h4925;
mem_array[8400] = 16'h3dc8;
mem_array[8403] = 16'haf1a;
mem_array[8402] = 16'hbda7;
mem_array[8405] = 16'h6a18;
mem_array[8404] = 16'hbd8f;
mem_array[8407] = 16'h9ae0;
mem_array[8406] = 16'h3cdc;
mem_array[8409] = 16'h6140;
mem_array[8408] = 16'hbd50;
mem_array[8411] = 16'h1a90;
mem_array[8410] = 16'hbd86;
mem_array[8413] = 16'he572;
mem_array[8412] = 16'h3c9c;
mem_array[8415] = 16'h9cd5;
mem_array[8414] = 16'h3d9d;
mem_array[8417] = 16'hbfc3;
mem_array[8416] = 16'hbd85;
mem_array[8419] = 16'hc129;
mem_array[8418] = 16'h3d24;
mem_array[8421] = 16'ha800;
mem_array[8420] = 16'h3c0c;
mem_array[8423] = 16'h5c2a;
mem_array[8422] = 16'h3d2c;
mem_array[8425] = 16'h1ee2;
mem_array[8424] = 16'hbd47;
mem_array[8427] = 16'h5c82;
mem_array[8426] = 16'hbdaa;
mem_array[8429] = 16'hc1d4;
mem_array[8428] = 16'h3d84;
mem_array[8431] = 16'h6c74;
mem_array[8430] = 16'h3bbf;
mem_array[8433] = 16'h2e62;
mem_array[8432] = 16'hbc9a;
mem_array[8435] = 16'hb0bd;
mem_array[8434] = 16'h3d52;
mem_array[8437] = 16'h52ae;
mem_array[8436] = 16'hbbba;
mem_array[8439] = 16'h74e6;
mem_array[8438] = 16'h3b82;
mem_array[8441] = 16'h84b6;
mem_array[8440] = 16'h3d90;
mem_array[8443] = 16'h1eea;
mem_array[8442] = 16'hbd46;
mem_array[8445] = 16'h5c6b;
mem_array[8444] = 16'h3b05;
mem_array[8447] = 16'h0583;
mem_array[8446] = 16'hbd5c;
mem_array[8449] = 16'h4c6f;
mem_array[8448] = 16'h3d8e;
mem_array[8451] = 16'h577f;
mem_array[8450] = 16'hbd87;
mem_array[8453] = 16'h2aaa;
mem_array[8452] = 16'hbd29;
mem_array[8455] = 16'h3a60;
mem_array[8454] = 16'hbda7;
mem_array[8457] = 16'he4cc;
mem_array[8456] = 16'h3d29;
mem_array[8459] = 16'h1907;
mem_array[8458] = 16'hbcd6;
mem_array[8461] = 16'h386c;
mem_array[8460] = 16'hba98;
mem_array[8463] = 16'he2fa;
mem_array[8462] = 16'hbb98;
mem_array[8465] = 16'h7dae;
mem_array[8464] = 16'h3d23;
mem_array[8467] = 16'h5938;
mem_array[8466] = 16'h3da4;
mem_array[8469] = 16'h61e5;
mem_array[8468] = 16'h3c48;
mem_array[8471] = 16'hfcbd;
mem_array[8470] = 16'h3dd0;
mem_array[8473] = 16'h4c95;
mem_array[8472] = 16'hbd75;
mem_array[8475] = 16'h2369;
mem_array[8474] = 16'h3d60;
mem_array[8477] = 16'h0219;
mem_array[8476] = 16'hbdd3;
mem_array[8479] = 16'h840b;
mem_array[8478] = 16'hbd5b;
mem_array[8481] = 16'h798b;
mem_array[8480] = 16'h3de0;
mem_array[8483] = 16'h007c;
mem_array[8482] = 16'hbad7;
mem_array[8485] = 16'h28ff;
mem_array[8484] = 16'hbc39;
mem_array[8487] = 16'h826c;
mem_array[8486] = 16'hbd74;
mem_array[8489] = 16'haf43;
mem_array[8488] = 16'h3d0a;
mem_array[8491] = 16'h1fc6;
mem_array[8490] = 16'h3dbd;
mem_array[8493] = 16'h6ab8;
mem_array[8492] = 16'h3da2;
mem_array[8495] = 16'h6f4a;
mem_array[8494] = 16'hbc9c;
mem_array[8497] = 16'h7031;
mem_array[8496] = 16'h3d61;
mem_array[8499] = 16'hce45;
mem_array[8498] = 16'hbdb5;
mem_array[8501] = 16'hf35d;
mem_array[8500] = 16'h3c9c;
mem_array[8503] = 16'h2211;
mem_array[8502] = 16'hbd9b;
mem_array[8505] = 16'h7e03;
mem_array[8504] = 16'h3db3;
mem_array[8507] = 16'h84b5;
mem_array[8506] = 16'hbdde;
mem_array[8509] = 16'h80d7;
mem_array[8508] = 16'hbd19;
mem_array[8511] = 16'h6657;
mem_array[8510] = 16'h3d9c;
mem_array[8513] = 16'h0ff5;
mem_array[8512] = 16'hbcc0;
mem_array[8515] = 16'h291a;
mem_array[8514] = 16'h3cd1;
mem_array[8517] = 16'h1846;
mem_array[8516] = 16'hbd30;
mem_array[8519] = 16'h27ee;
mem_array[8518] = 16'hbd08;
mem_array[8521] = 16'h953d;
mem_array[8520] = 16'h3ee2;
mem_array[8523] = 16'h421f;
mem_array[8522] = 16'hbde1;
mem_array[8525] = 16'h1272;
mem_array[8524] = 16'h3ef5;
mem_array[8527] = 16'hc144;
mem_array[8526] = 16'hbe29;
mem_array[8529] = 16'h2c2e;
mem_array[8528] = 16'h3c90;
mem_array[8531] = 16'h9e38;
mem_array[8530] = 16'h3cca;
mem_array[8533] = 16'hcd26;
mem_array[8532] = 16'h3e90;
mem_array[8535] = 16'h864c;
mem_array[8534] = 16'h3e83;
mem_array[8537] = 16'h8b85;
mem_array[8536] = 16'hbdc0;
mem_array[8539] = 16'hf8e5;
mem_array[8538] = 16'h3f4f;
mem_array[8541] = 16'hc427;
mem_array[8540] = 16'h3ce9;
mem_array[8543] = 16'h8243;
mem_array[8542] = 16'hbd17;
mem_array[8545] = 16'h9738;
mem_array[8544] = 16'hbe93;
mem_array[8547] = 16'h8c90;
mem_array[8546] = 16'h3f46;
mem_array[8549] = 16'h3666;
mem_array[8548] = 16'h3ed7;
mem_array[8551] = 16'h6519;
mem_array[8550] = 16'h3f69;
mem_array[8553] = 16'h776f;
mem_array[8552] = 16'h3e39;
mem_array[8555] = 16'h05c0;
mem_array[8554] = 16'hbdbe;
mem_array[8557] = 16'h72c3;
mem_array[8556] = 16'h3c81;
mem_array[8559] = 16'h835e;
mem_array[8558] = 16'h3cb8;
mem_array[8561] = 16'hf1b7;
mem_array[8560] = 16'hbe8a;
mem_array[8563] = 16'h55e3;
mem_array[8562] = 16'hbe04;
mem_array[8565] = 16'hd9b1;
mem_array[8564] = 16'hbf38;
mem_array[8567] = 16'h8f91;
mem_array[8566] = 16'hbf7b;
mem_array[8569] = 16'hd945;
mem_array[8568] = 16'h3edd;
mem_array[8571] = 16'h399a;
mem_array[8570] = 16'hbd50;
mem_array[8573] = 16'h49bd;
mem_array[8572] = 16'h3e5e;
mem_array[8575] = 16'h50c6;
mem_array[8574] = 16'hbd7b;
mem_array[8577] = 16'h595e;
mem_array[8576] = 16'hbc18;
mem_array[8579] = 16'h6433;
mem_array[8578] = 16'hbed9;
mem_array[8581] = 16'h96b3;
mem_array[8580] = 16'h3f4a;
mem_array[8583] = 16'h102a;
mem_array[8582] = 16'hbe58;
mem_array[8585] = 16'h2a20;
mem_array[8584] = 16'hbe9e;
mem_array[8587] = 16'hf666;
mem_array[8586] = 16'h3e5b;
mem_array[8589] = 16'h9dd6;
mem_array[8588] = 16'h3e62;
mem_array[8591] = 16'h035d;
mem_array[8590] = 16'h3cc4;
mem_array[8593] = 16'h309f;
mem_array[8592] = 16'h3f16;
mem_array[8595] = 16'h1036;
mem_array[8594] = 16'h3e75;
mem_array[8597] = 16'h1dd9;
mem_array[8596] = 16'hbe79;
mem_array[8599] = 16'hae7a;
mem_array[8598] = 16'h3f1a;
mem_array[8601] = 16'h2025;
mem_array[8600] = 16'h3ca1;
mem_array[8603] = 16'h422e;
mem_array[8602] = 16'h3d9e;
mem_array[8605] = 16'heec0;
mem_array[8604] = 16'h3e2c;
mem_array[8607] = 16'hd84d;
mem_array[8606] = 16'h3e10;
mem_array[8609] = 16'h0c93;
mem_array[8608] = 16'h3d9b;
mem_array[8611] = 16'h6fee;
mem_array[8610] = 16'hbd8e;
mem_array[8613] = 16'hb559;
mem_array[8612] = 16'h3e99;
mem_array[8615] = 16'h8d41;
mem_array[8614] = 16'h3cee;
mem_array[8617] = 16'h7599;
mem_array[8616] = 16'h3e6d;
mem_array[8619] = 16'h6539;
mem_array[8618] = 16'h3bf5;
mem_array[8621] = 16'hc054;
mem_array[8620] = 16'hbe55;
mem_array[8623] = 16'h527c;
mem_array[8622] = 16'h3c62;
mem_array[8625] = 16'hb886;
mem_array[8624] = 16'hbf1d;
mem_array[8627] = 16'h7319;
mem_array[8626] = 16'hbe6f;
mem_array[8629] = 16'h4551;
mem_array[8628] = 16'h3f6c;
mem_array[8631] = 16'h397e;
mem_array[8630] = 16'h3f17;
mem_array[8633] = 16'h67d1;
mem_array[8632] = 16'h3f74;
mem_array[8635] = 16'hf0d7;
mem_array[8634] = 16'h3e02;
mem_array[8637] = 16'h474d;
mem_array[8636] = 16'hbe7d;
mem_array[8639] = 16'h07ba;
mem_array[8638] = 16'hbf5f;
mem_array[8641] = 16'he5bc;
mem_array[8640] = 16'hbd8f;
mem_array[8643] = 16'ha205;
mem_array[8642] = 16'hbecc;
mem_array[8645] = 16'hf189;
mem_array[8644] = 16'h3f22;
mem_array[8647] = 16'h3e6c;
mem_array[8646] = 16'h3f4c;
mem_array[8649] = 16'hc942;
mem_array[8648] = 16'h3ed4;
mem_array[8651] = 16'hfda1;
mem_array[8650] = 16'hbf04;
mem_array[8653] = 16'h2356;
mem_array[8652] = 16'h3f84;
mem_array[8655] = 16'hee04;
mem_array[8654] = 16'h3edc;
mem_array[8657] = 16'h5752;
mem_array[8656] = 16'h3d40;
mem_array[8659] = 16'hf1d8;
mem_array[8658] = 16'hbf5b;
mem_array[8661] = 16'hf79e;
mem_array[8660] = 16'hbdb9;
mem_array[8663] = 16'hd3f7;
mem_array[8662] = 16'hbbbd;
mem_array[8665] = 16'hb3a4;
mem_array[8664] = 16'hbf62;
mem_array[8667] = 16'h6cf4;
mem_array[8666] = 16'h3f0d;
mem_array[8669] = 16'hc059;
mem_array[8668] = 16'h3ee7;
mem_array[8671] = 16'h8d26;
mem_array[8670] = 16'hbef7;
mem_array[8673] = 16'h2e77;
mem_array[8672] = 16'h3ec3;
mem_array[8675] = 16'h2da4;
mem_array[8674] = 16'h3e06;
mem_array[8677] = 16'h26c4;
mem_array[8676] = 16'hbfba;
mem_array[8679] = 16'h9248;
mem_array[8678] = 16'h3e1f;
mem_array[8681] = 16'h72eb;
mem_array[8680] = 16'hbd2e;
mem_array[8683] = 16'hd209;
mem_array[8682] = 16'h3e6e;
mem_array[8685] = 16'hb5bd;
mem_array[8684] = 16'hbdbf;
mem_array[8687] = 16'h0ccd;
mem_array[8686] = 16'h3ef1;
mem_array[8689] = 16'hf13c;
mem_array[8688] = 16'hbd10;
mem_array[8691] = 16'hf796;
mem_array[8690] = 16'hbec6;
mem_array[8693] = 16'h57ab;
mem_array[8692] = 16'h3dea;
mem_array[8695] = 16'h53bf;
mem_array[8694] = 16'h3f2f;
mem_array[8697] = 16'h0fda;
mem_array[8696] = 16'h3bb4;
mem_array[8699] = 16'h127d;
mem_array[8698] = 16'hbc67;
mem_array[8701] = 16'h1a76;
mem_array[8700] = 16'h3e91;
mem_array[8703] = 16'h1d46;
mem_array[8702] = 16'hbf14;
mem_array[8705] = 16'hb376;
mem_array[8704] = 16'hbf8c;
mem_array[8707] = 16'h64ba;
mem_array[8706] = 16'hbf45;
mem_array[8709] = 16'hdd10;
mem_array[8708] = 16'h3dad;
mem_array[8711] = 16'h6e47;
mem_array[8710] = 16'hbfab;
mem_array[8713] = 16'h8be8;
mem_array[8712] = 16'h3f5a;
mem_array[8715] = 16'hb23e;
mem_array[8714] = 16'hbed2;
mem_array[8717] = 16'h176f;
mem_array[8716] = 16'hbe5f;
mem_array[8719] = 16'h09ce;
mem_array[8718] = 16'h3e7d;
mem_array[8721] = 16'h0a73;
mem_array[8720] = 16'h3d70;
mem_array[8723] = 16'h7812;
mem_array[8722] = 16'hbd58;
mem_array[8725] = 16'hdcbf;
mem_array[8724] = 16'hbf08;
mem_array[8727] = 16'h7f07;
mem_array[8726] = 16'hbf04;
mem_array[8729] = 16'h7456;
mem_array[8728] = 16'h3e94;
mem_array[8731] = 16'h20c6;
mem_array[8730] = 16'h3e52;
mem_array[8733] = 16'h1e01;
mem_array[8732] = 16'hbed0;
mem_array[8735] = 16'hc7cd;
mem_array[8734] = 16'h3e14;
mem_array[8737] = 16'hae68;
mem_array[8736] = 16'hbf10;
mem_array[8739] = 16'hb508;
mem_array[8738] = 16'h3d96;
mem_array[8741] = 16'h2de1;
mem_array[8740] = 16'hbea7;
mem_array[8743] = 16'h2a5e;
mem_array[8742] = 16'h3e80;
mem_array[8745] = 16'h8fc8;
mem_array[8744] = 16'hbf24;
mem_array[8747] = 16'hde7a;
mem_array[8746] = 16'h3e58;
mem_array[8749] = 16'h5ef1;
mem_array[8748] = 16'hbea2;
mem_array[8751] = 16'h00a9;
mem_array[8750] = 16'h3d83;
mem_array[8753] = 16'hca98;
mem_array[8752] = 16'hbea7;
mem_array[8755] = 16'h6536;
mem_array[8754] = 16'h3ecb;
mem_array[8757] = 16'h6391;
mem_array[8756] = 16'hbe95;
mem_array[8759] = 16'h77a0;
mem_array[8758] = 16'hbe68;
mem_array[8761] = 16'hc00d;
mem_array[8760] = 16'hbe8b;
mem_array[8763] = 16'h54c6;
mem_array[8762] = 16'hbfbe;
mem_array[8765] = 16'h4bbe;
mem_array[8764] = 16'hbf18;
mem_array[8767] = 16'hc962;
mem_array[8766] = 16'hbe33;
mem_array[8769] = 16'h84d9;
mem_array[8768] = 16'h3e8a;
mem_array[8771] = 16'h2e2b;
mem_array[8770] = 16'hbf8c;
mem_array[8773] = 16'hf761;
mem_array[8772] = 16'h3f04;
mem_array[8775] = 16'h966a;
mem_array[8774] = 16'h3d31;
mem_array[8777] = 16'h66fb;
mem_array[8776] = 16'h3eb7;
mem_array[8779] = 16'hcdef;
mem_array[8778] = 16'h3ea4;
mem_array[8781] = 16'h78fa;
mem_array[8780] = 16'hba93;
mem_array[8783] = 16'h8d2f;
mem_array[8782] = 16'hbd0a;
mem_array[8785] = 16'h1947;
mem_array[8784] = 16'h3eb6;
mem_array[8787] = 16'hb252;
mem_array[8786] = 16'h3e98;
mem_array[8789] = 16'h201b;
mem_array[8788] = 16'h3db6;
mem_array[8791] = 16'h3e0e;
mem_array[8790] = 16'hbda3;
mem_array[8793] = 16'hfa97;
mem_array[8792] = 16'hbe2b;
mem_array[8795] = 16'h1a2c;
mem_array[8794] = 16'h3dc4;
mem_array[8797] = 16'hc8c3;
mem_array[8796] = 16'hbf81;
mem_array[8799] = 16'hc05e;
mem_array[8798] = 16'h3e25;
mem_array[8801] = 16'hece7;
mem_array[8800] = 16'h3d7d;
mem_array[8803] = 16'haecf;
mem_array[8802] = 16'h3edc;
mem_array[8805] = 16'hfc16;
mem_array[8804] = 16'hbf8b;
mem_array[8807] = 16'h70a3;
mem_array[8806] = 16'h3e28;
mem_array[8809] = 16'h8eb3;
mem_array[8808] = 16'hbec9;
mem_array[8811] = 16'h8b49;
mem_array[8810] = 16'hbf17;
mem_array[8813] = 16'hd0ca;
mem_array[8812] = 16'hbf19;
mem_array[8815] = 16'ha3a7;
mem_array[8814] = 16'h3e38;
mem_array[8817] = 16'h1e3d;
mem_array[8816] = 16'h3d87;
mem_array[8819] = 16'h7907;
mem_array[8818] = 16'hbf58;
mem_array[8821] = 16'he197;
mem_array[8820] = 16'hbe53;
mem_array[8823] = 16'hb4e7;
mem_array[8822] = 16'hbfb9;
mem_array[8825] = 16'h4516;
mem_array[8824] = 16'h3ed0;
mem_array[8827] = 16'h1c4e;
mem_array[8826] = 16'hbe6e;
mem_array[8829] = 16'h2f52;
mem_array[8828] = 16'h3f3d;
mem_array[8831] = 16'h44c0;
mem_array[8830] = 16'hbe1c;
mem_array[8833] = 16'hf566;
mem_array[8832] = 16'h3e5d;
mem_array[8835] = 16'hcf02;
mem_array[8834] = 16'h3e1c;
mem_array[8837] = 16'h1d76;
mem_array[8836] = 16'h3e89;
mem_array[8839] = 16'h5d45;
mem_array[8838] = 16'hbe14;
mem_array[8841] = 16'h14ec;
mem_array[8840] = 16'h3a28;
mem_array[8843] = 16'h6d7b;
mem_array[8842] = 16'h3dae;
mem_array[8845] = 16'hea14;
mem_array[8844] = 16'h3cf1;
mem_array[8847] = 16'h6fa3;
mem_array[8846] = 16'h3e8b;
mem_array[8849] = 16'h8f23;
mem_array[8848] = 16'hbe97;
mem_array[8851] = 16'he884;
mem_array[8850] = 16'hbe92;
mem_array[8853] = 16'h3e1d;
mem_array[8852] = 16'h3ec9;
mem_array[8855] = 16'h1c7f;
mem_array[8854] = 16'h3cc8;
mem_array[8857] = 16'hae7e;
mem_array[8856] = 16'h3dc6;
mem_array[8859] = 16'h3516;
mem_array[8858] = 16'hbcea;
mem_array[8861] = 16'haf77;
mem_array[8860] = 16'h3ef4;
mem_array[8863] = 16'h8e85;
mem_array[8862] = 16'h3e6b;
mem_array[8865] = 16'h3940;
mem_array[8864] = 16'hbfbe;
mem_array[8867] = 16'h6f44;
mem_array[8866] = 16'h3f08;
mem_array[8869] = 16'h8462;
mem_array[8868] = 16'hbd9e;
mem_array[8871] = 16'h18b4;
mem_array[8870] = 16'h3d55;
mem_array[8873] = 16'hef9c;
mem_array[8872] = 16'hbf22;
mem_array[8875] = 16'h8a74;
mem_array[8874] = 16'hbdf8;
mem_array[8877] = 16'h297c;
mem_array[8876] = 16'hbe38;
mem_array[8879] = 16'hd70c;
mem_array[8878] = 16'hbf3d;
mem_array[8881] = 16'h59df;
mem_array[8880] = 16'hbfc4;
mem_array[8883] = 16'h63bf;
mem_array[8882] = 16'hbdcd;
mem_array[8885] = 16'hf8c9;
mem_array[8884] = 16'h3e4c;
mem_array[8887] = 16'hcf60;
mem_array[8886] = 16'hbe4b;
mem_array[8889] = 16'h8eb4;
mem_array[8888] = 16'h3f86;
mem_array[8891] = 16'h4040;
mem_array[8890] = 16'hbc67;
mem_array[8893] = 16'h5e47;
mem_array[8892] = 16'h3cb2;
mem_array[8895] = 16'h4f11;
mem_array[8894] = 16'h3db9;
mem_array[8897] = 16'h5260;
mem_array[8896] = 16'hbe03;
mem_array[8899] = 16'hea09;
mem_array[8898] = 16'hbf46;
mem_array[8901] = 16'h6cbf;
mem_array[8900] = 16'h3d71;
mem_array[8903] = 16'h35ef;
mem_array[8902] = 16'hbd6c;
mem_array[8905] = 16'h2f4e;
mem_array[8904] = 16'hbd27;
mem_array[8907] = 16'h94bf;
mem_array[8906] = 16'hbc58;
mem_array[8909] = 16'h164b;
mem_array[8908] = 16'hbeda;
mem_array[8911] = 16'hd68c;
mem_array[8910] = 16'hbdfa;
mem_array[8913] = 16'hbf95;
mem_array[8912] = 16'h3d9c;
mem_array[8915] = 16'hc79e;
mem_array[8914] = 16'hbef2;
mem_array[8917] = 16'h45f2;
mem_array[8916] = 16'h3f0b;
mem_array[8919] = 16'hbfad;
mem_array[8918] = 16'hbe7a;
mem_array[8921] = 16'heb84;
mem_array[8920] = 16'h3e5f;
mem_array[8923] = 16'hf995;
mem_array[8922] = 16'h3ef4;
mem_array[8925] = 16'hed8e;
mem_array[8924] = 16'h3f34;
mem_array[8927] = 16'hc784;
mem_array[8926] = 16'h3e34;
mem_array[8929] = 16'h071a;
mem_array[8928] = 16'hbe3f;
mem_array[8931] = 16'hf566;
mem_array[8930] = 16'h3f51;
mem_array[8933] = 16'h5f0f;
mem_array[8932] = 16'hbe2a;
mem_array[8935] = 16'h32a0;
mem_array[8934] = 16'h3d0f;
mem_array[8937] = 16'h7433;
mem_array[8936] = 16'hbe85;
mem_array[8939] = 16'ha7fe;
mem_array[8938] = 16'hbf00;
mem_array[8941] = 16'hebf6;
mem_array[8940] = 16'h3db5;
mem_array[8943] = 16'h13d8;
mem_array[8942] = 16'hbdaa;
mem_array[8945] = 16'h66b2;
mem_array[8944] = 16'h3e89;
mem_array[8947] = 16'h5b43;
mem_array[8946] = 16'hbe64;
mem_array[8949] = 16'h2c31;
mem_array[8948] = 16'h3f3a;
mem_array[8951] = 16'h66d8;
mem_array[8950] = 16'hbe4c;
mem_array[8953] = 16'h69ed;
mem_array[8952] = 16'hbde2;
mem_array[8955] = 16'h7d98;
mem_array[8954] = 16'h3ecb;
mem_array[8957] = 16'ha959;
mem_array[8956] = 16'hbeaf;
mem_array[8959] = 16'h3495;
mem_array[8958] = 16'hbf15;
mem_array[8961] = 16'hc0fc;
mem_array[8960] = 16'hbd56;
mem_array[8963] = 16'h2ec2;
mem_array[8962] = 16'h3d95;
mem_array[8965] = 16'he14f;
mem_array[8964] = 16'h3df1;
mem_array[8967] = 16'hd5ea;
mem_array[8966] = 16'h3e77;
mem_array[8969] = 16'hc742;
mem_array[8968] = 16'hbf21;
mem_array[8971] = 16'h9fd1;
mem_array[8970] = 16'hbdfd;
mem_array[8973] = 16'hb151;
mem_array[8972] = 16'h3e13;
mem_array[8975] = 16'h3c07;
mem_array[8974] = 16'hbdd2;
mem_array[8977] = 16'hdd53;
mem_array[8976] = 16'hbeb3;
mem_array[8979] = 16'ha150;
mem_array[8978] = 16'h3dc3;
mem_array[8981] = 16'hfed1;
mem_array[8980] = 16'hbe81;
mem_array[8983] = 16'h7849;
mem_array[8982] = 16'h3e81;
mem_array[8985] = 16'hdcea;
mem_array[8984] = 16'h3e81;
mem_array[8987] = 16'h60de;
mem_array[8986] = 16'h3e68;
mem_array[8989] = 16'h0f12;
mem_array[8988] = 16'hbe90;
mem_array[8991] = 16'h07a7;
mem_array[8990] = 16'h3ef2;
mem_array[8993] = 16'he41e;
mem_array[8992] = 16'h3ca4;
mem_array[8995] = 16'h3e74;
mem_array[8994] = 16'hbef3;
mem_array[8997] = 16'h16d2;
mem_array[8996] = 16'h3db9;
mem_array[8999] = 16'h1a91;
mem_array[8998] = 16'hbec0;
mem_array[9001] = 16'h87ab;
mem_array[9000] = 16'hbfd9;
mem_array[9003] = 16'h398d;
mem_array[9002] = 16'hbfa1;
mem_array[9005] = 16'hed34;
mem_array[9004] = 16'h3e35;
mem_array[9007] = 16'h4c22;
mem_array[9006] = 16'hbe3c;
mem_array[9009] = 16'hf24b;
mem_array[9008] = 16'h3ea3;
mem_array[9011] = 16'hecf1;
mem_array[9010] = 16'h3ee7;
mem_array[9013] = 16'h39af;
mem_array[9012] = 16'h3d10;
mem_array[9015] = 16'h476d;
mem_array[9014] = 16'h3e47;
mem_array[9017] = 16'h54e8;
mem_array[9016] = 16'hbe2e;
mem_array[9019] = 16'hf2f8;
mem_array[9018] = 16'hbef4;
mem_array[9021] = 16'h3819;
mem_array[9020] = 16'hbd90;
mem_array[9023] = 16'h41a4;
mem_array[9022] = 16'hbd3e;
mem_array[9025] = 16'hf0de;
mem_array[9024] = 16'h3eb9;
mem_array[9027] = 16'hd5ae;
mem_array[9026] = 16'h3e63;
mem_array[9029] = 16'h2d78;
mem_array[9028] = 16'hbe91;
mem_array[9031] = 16'h83e6;
mem_array[9030] = 16'hbda7;
mem_array[9033] = 16'hebc3;
mem_array[9032] = 16'hbec3;
mem_array[9035] = 16'h224d;
mem_array[9034] = 16'h3e5c;
mem_array[9037] = 16'ha656;
mem_array[9036] = 16'hbe8c;
mem_array[9039] = 16'h437d;
mem_array[9038] = 16'h3c94;
mem_array[9041] = 16'hb539;
mem_array[9040] = 16'hbe25;
mem_array[9043] = 16'h71ed;
mem_array[9042] = 16'hbd5d;
mem_array[9045] = 16'h096c;
mem_array[9044] = 16'hbdf3;
mem_array[9047] = 16'h674e;
mem_array[9046] = 16'hbe8b;
mem_array[9049] = 16'ha3c8;
mem_array[9048] = 16'hbe91;
mem_array[9051] = 16'hb51d;
mem_array[9050] = 16'hbeb4;
mem_array[9053] = 16'h973c;
mem_array[9052] = 16'hbe64;
mem_array[9055] = 16'h4985;
mem_array[9054] = 16'hbcac;
mem_array[9057] = 16'h0004;
mem_array[9056] = 16'h3e24;
mem_array[9059] = 16'ha7dc;
mem_array[9058] = 16'hbe3e;
mem_array[9061] = 16'h99c1;
mem_array[9060] = 16'hbfd8;
mem_array[9063] = 16'h19c6;
mem_array[9062] = 16'hbe6c;
mem_array[9065] = 16'hbe6f;
mem_array[9064] = 16'hbc83;
mem_array[9067] = 16'hed95;
mem_array[9066] = 16'hbe46;
mem_array[9069] = 16'h1679;
mem_array[9068] = 16'hbe30;
mem_array[9071] = 16'h28b3;
mem_array[9070] = 16'h3d87;
mem_array[9073] = 16'hf21f;
mem_array[9072] = 16'h3dd2;
mem_array[9075] = 16'hb3fb;
mem_array[9074] = 16'h3d80;
mem_array[9077] = 16'h6c0d;
mem_array[9076] = 16'h3e80;
mem_array[9079] = 16'hf343;
mem_array[9078] = 16'hbd8c;
mem_array[9081] = 16'hb339;
mem_array[9080] = 16'hbcc1;
mem_array[9083] = 16'hd1af;
mem_array[9082] = 16'h3cfc;
mem_array[9085] = 16'hd396;
mem_array[9084] = 16'hbe58;
mem_array[9087] = 16'ha114;
mem_array[9086] = 16'h3e0c;
mem_array[9089] = 16'h41ed;
mem_array[9088] = 16'hbea5;
mem_array[9091] = 16'h5696;
mem_array[9090] = 16'h3db6;
mem_array[9093] = 16'h6bc5;
mem_array[9092] = 16'h3db7;
mem_array[9095] = 16'h0e08;
mem_array[9094] = 16'hbc71;
mem_array[9097] = 16'h9c40;
mem_array[9096] = 16'hbd11;
mem_array[9099] = 16'h0b72;
mem_array[9098] = 16'hbdad;
mem_array[9101] = 16'h4e7f;
mem_array[9100] = 16'hbd6b;
mem_array[9103] = 16'h7087;
mem_array[9102] = 16'h3d9f;
mem_array[9105] = 16'h2fb7;
mem_array[9104] = 16'hbe4c;
mem_array[9107] = 16'h178f;
mem_array[9106] = 16'hbd99;
mem_array[9109] = 16'h55f6;
mem_array[9108] = 16'h3d86;
mem_array[9111] = 16'h3148;
mem_array[9110] = 16'hbe63;
mem_array[9113] = 16'hf3cf;
mem_array[9112] = 16'h3e3c;
mem_array[9115] = 16'hba1b;
mem_array[9114] = 16'hbdaa;
mem_array[9117] = 16'h0ea1;
mem_array[9116] = 16'h3e51;
mem_array[9119] = 16'hfee6;
mem_array[9118] = 16'hbebd;
mem_array[9121] = 16'h6871;
mem_array[9120] = 16'hbf6d;
mem_array[9123] = 16'h7933;
mem_array[9122] = 16'h3c34;
mem_array[9125] = 16'h8c4b;
mem_array[9124] = 16'h3e7b;
mem_array[9127] = 16'h7da1;
mem_array[9126] = 16'hbcd3;
mem_array[9129] = 16'hc403;
mem_array[9128] = 16'h3dfe;
mem_array[9131] = 16'he353;
mem_array[9130] = 16'hbd43;
mem_array[9133] = 16'h38c8;
mem_array[9132] = 16'h3dc5;
mem_array[9135] = 16'h6241;
mem_array[9134] = 16'h3ee8;
mem_array[9137] = 16'hb391;
mem_array[9136] = 16'h3e5d;
mem_array[9139] = 16'hf3eb;
mem_array[9138] = 16'hbdad;
mem_array[9141] = 16'he3de;
mem_array[9140] = 16'h3c80;
mem_array[9143] = 16'h8dd1;
mem_array[9142] = 16'hbd0f;
mem_array[9145] = 16'h3245;
mem_array[9144] = 16'h3d99;
mem_array[9147] = 16'ha4b4;
mem_array[9146] = 16'h3e5b;
mem_array[9149] = 16'h5956;
mem_array[9148] = 16'hbe7c;
mem_array[9151] = 16'h520d;
mem_array[9150] = 16'hbdd3;
mem_array[9153] = 16'h3c8a;
mem_array[9152] = 16'h3e8c;
mem_array[9155] = 16'h7b17;
mem_array[9154] = 16'hbc91;
mem_array[9157] = 16'h84cf;
mem_array[9156] = 16'h3e3f;
mem_array[9159] = 16'h49d2;
mem_array[9158] = 16'hbe9e;
mem_array[9161] = 16'hc34e;
mem_array[9160] = 16'h3d3d;
mem_array[9163] = 16'h6a35;
mem_array[9162] = 16'hbccb;
mem_array[9165] = 16'hff95;
mem_array[9164] = 16'hbdaf;
mem_array[9167] = 16'h5927;
mem_array[9166] = 16'h3def;
mem_array[9169] = 16'h4e99;
mem_array[9168] = 16'hbe53;
mem_array[9171] = 16'hb923;
mem_array[9170] = 16'h3df2;
mem_array[9173] = 16'h48b2;
mem_array[9172] = 16'hbda5;
mem_array[9175] = 16'h7e3d;
mem_array[9174] = 16'hbe21;
mem_array[9177] = 16'h9303;
mem_array[9176] = 16'h3d1a;
mem_array[9179] = 16'h0cbe;
mem_array[9178] = 16'hbf45;
mem_array[9181] = 16'h8ceb;
mem_array[9180] = 16'hbf80;
mem_array[9183] = 16'hcd7b;
mem_array[9182] = 16'hbf10;
mem_array[9185] = 16'h074a;
mem_array[9184] = 16'h3df4;
mem_array[9187] = 16'h512d;
mem_array[9186] = 16'hbd51;
mem_array[9189] = 16'h09d4;
mem_array[9188] = 16'hbdc1;
mem_array[9191] = 16'hae92;
mem_array[9190] = 16'hbdab;
mem_array[9193] = 16'h5ec3;
mem_array[9192] = 16'h3e66;
mem_array[9195] = 16'hddd5;
mem_array[9194] = 16'h3ea2;
mem_array[9197] = 16'h1292;
mem_array[9196] = 16'hbb9c;
mem_array[9199] = 16'hdd72;
mem_array[9198] = 16'hbe6c;
mem_array[9201] = 16'hc834;
mem_array[9200] = 16'h3d77;
mem_array[9203] = 16'hf47b;
mem_array[9202] = 16'hbdb3;
mem_array[9205] = 16'h7641;
mem_array[9204] = 16'h3e6c;
mem_array[9207] = 16'hc459;
mem_array[9206] = 16'h3eae;
mem_array[9209] = 16'h1e6a;
mem_array[9208] = 16'hbe17;
mem_array[9211] = 16'hb44e;
mem_array[9210] = 16'hbde2;
mem_array[9213] = 16'h3181;
mem_array[9212] = 16'h3e60;
mem_array[9215] = 16'hf52f;
mem_array[9214] = 16'hbdec;
mem_array[9217] = 16'heb97;
mem_array[9216] = 16'hbeb3;
mem_array[9219] = 16'h4aeb;
mem_array[9218] = 16'hbea3;
mem_array[9221] = 16'he48a;
mem_array[9220] = 16'h3e30;
mem_array[9223] = 16'hbdc2;
mem_array[9222] = 16'hbe15;
mem_array[9225] = 16'hde2d;
mem_array[9224] = 16'hbe92;
mem_array[9227] = 16'h9bd7;
mem_array[9226] = 16'h3e35;
mem_array[9229] = 16'h28e9;
mem_array[9228] = 16'h3c30;
mem_array[9231] = 16'h41f1;
mem_array[9230] = 16'hbedc;
mem_array[9233] = 16'h0166;
mem_array[9232] = 16'hbe7d;
mem_array[9235] = 16'hf099;
mem_array[9234] = 16'hbe08;
mem_array[9237] = 16'hf6b2;
mem_array[9236] = 16'h3d4f;
mem_array[9239] = 16'h8978;
mem_array[9238] = 16'hbec7;
mem_array[9241] = 16'h8d35;
mem_array[9240] = 16'hbed8;
mem_array[9243] = 16'h924a;
mem_array[9242] = 16'hbe99;
mem_array[9245] = 16'h8128;
mem_array[9244] = 16'hbe3b;
mem_array[9247] = 16'h901f;
mem_array[9246] = 16'h3cce;
mem_array[9249] = 16'h48c2;
mem_array[9248] = 16'hbd23;
mem_array[9251] = 16'h8c76;
mem_array[9250] = 16'hba8d;
mem_array[9253] = 16'hdd5a;
mem_array[9252] = 16'hbd87;
mem_array[9255] = 16'h918c;
mem_array[9254] = 16'h3dc7;
mem_array[9257] = 16'hb186;
mem_array[9256] = 16'hbec9;
mem_array[9259] = 16'h07ee;
mem_array[9258] = 16'hbd8b;
mem_array[9261] = 16'h8b7f;
mem_array[9260] = 16'hbdca;
mem_array[9263] = 16'h15de;
mem_array[9262] = 16'h3c98;
mem_array[9265] = 16'h2ff2;
mem_array[9264] = 16'hbe2a;
mem_array[9267] = 16'hc744;
mem_array[9266] = 16'h3e99;
mem_array[9269] = 16'hf182;
mem_array[9268] = 16'hbeaa;
mem_array[9271] = 16'h10e0;
mem_array[9270] = 16'h3d50;
mem_array[9273] = 16'h1455;
mem_array[9272] = 16'hbdbc;
mem_array[9275] = 16'h155c;
mem_array[9274] = 16'hbf90;
mem_array[9277] = 16'h3648;
mem_array[9276] = 16'hbe81;
mem_array[9279] = 16'h1ec8;
mem_array[9278] = 16'h3dff;
mem_array[9281] = 16'hb4fe;
mem_array[9280] = 16'hbd24;
mem_array[9283] = 16'h5cc7;
mem_array[9282] = 16'hbcd5;
mem_array[9285] = 16'h1ef8;
mem_array[9284] = 16'hbe78;
mem_array[9287] = 16'h9fa8;
mem_array[9286] = 16'h3daa;
mem_array[9289] = 16'h8a9f;
mem_array[9288] = 16'hbda8;
mem_array[9291] = 16'h3e89;
mem_array[9290] = 16'hbee8;
mem_array[9293] = 16'haffc;
mem_array[9292] = 16'hbcf1;
mem_array[9295] = 16'h0132;
mem_array[9294] = 16'hbced;
mem_array[9297] = 16'h92bf;
mem_array[9296] = 16'h3e98;
mem_array[9299] = 16'h5426;
mem_array[9298] = 16'h3e6e;
mem_array[9301] = 16'h3646;
mem_array[9300] = 16'h3e8b;
mem_array[9303] = 16'h9b30;
mem_array[9302] = 16'hbf6e;
mem_array[9305] = 16'h694c;
mem_array[9304] = 16'hbd85;
mem_array[9307] = 16'h93af;
mem_array[9306] = 16'h3d88;
mem_array[9309] = 16'h2689;
mem_array[9308] = 16'hbe40;
mem_array[9311] = 16'h9004;
mem_array[9310] = 16'hbd81;
mem_array[9313] = 16'hd238;
mem_array[9312] = 16'h3e35;
mem_array[9315] = 16'h4e41;
mem_array[9314] = 16'h3e8a;
mem_array[9317] = 16'h3b56;
mem_array[9316] = 16'hbe9f;
mem_array[9319] = 16'h71b1;
mem_array[9318] = 16'h3e76;
mem_array[9321] = 16'h966f;
mem_array[9320] = 16'hbe19;
mem_array[9323] = 16'hd55c;
mem_array[9322] = 16'hbb84;
mem_array[9325] = 16'h0e33;
mem_array[9324] = 16'hbf00;
mem_array[9327] = 16'h954e;
mem_array[9326] = 16'h3e79;
mem_array[9329] = 16'h9ebf;
mem_array[9328] = 16'hbeac;
mem_array[9331] = 16'hb99a;
mem_array[9330] = 16'hbcf6;
mem_array[9333] = 16'hfe6b;
mem_array[9332] = 16'hbed5;
mem_array[9335] = 16'h26e5;
mem_array[9334] = 16'hbf55;
mem_array[9337] = 16'h47f7;
mem_array[9336] = 16'hbd72;
mem_array[9339] = 16'h4de6;
mem_array[9338] = 16'hbe72;
mem_array[9341] = 16'h24d8;
mem_array[9340] = 16'hbeaa;
mem_array[9343] = 16'h106a;
mem_array[9342] = 16'hbd76;
mem_array[9345] = 16'ha8fd;
mem_array[9344] = 16'hbe9f;
mem_array[9347] = 16'h29f2;
mem_array[9346] = 16'h3c36;
mem_array[9349] = 16'h1446;
mem_array[9348] = 16'hbd8e;
mem_array[9351] = 16'hf07e;
mem_array[9350] = 16'hbe8b;
mem_array[9353] = 16'h6445;
mem_array[9352] = 16'hbeb1;
mem_array[9355] = 16'h247c;
mem_array[9354] = 16'hbf04;
mem_array[9357] = 16'h9594;
mem_array[9356] = 16'h3e09;
mem_array[9359] = 16'hea52;
mem_array[9358] = 16'h3e60;
mem_array[9361] = 16'h5013;
mem_array[9360] = 16'hbdfc;
mem_array[9363] = 16'h30f5;
mem_array[9362] = 16'hbf2e;
mem_array[9365] = 16'h6708;
mem_array[9364] = 16'h3e05;
mem_array[9367] = 16'hea98;
mem_array[9366] = 16'h3e2e;
mem_array[9369] = 16'h9be1;
mem_array[9368] = 16'hbf07;
mem_array[9371] = 16'h933e;
mem_array[9370] = 16'hbb9e;
mem_array[9373] = 16'h5270;
mem_array[9372] = 16'hbd53;
mem_array[9375] = 16'h69f7;
mem_array[9374] = 16'h3e82;
mem_array[9377] = 16'h491e;
mem_array[9376] = 16'hbcfa;
mem_array[9379] = 16'h4c65;
mem_array[9378] = 16'h3e6c;
mem_array[9381] = 16'h71e0;
mem_array[9380] = 16'h3d3d;
mem_array[9383] = 16'hd4c2;
mem_array[9382] = 16'hbb06;
mem_array[9385] = 16'h4b1d;
mem_array[9384] = 16'hbf00;
mem_array[9387] = 16'h318f;
mem_array[9386] = 16'h3e9b;
mem_array[9389] = 16'hdb33;
mem_array[9388] = 16'h3e36;
mem_array[9391] = 16'h3112;
mem_array[9390] = 16'hbdbc;
mem_array[9393] = 16'h4ab5;
mem_array[9392] = 16'hbe7b;
mem_array[9395] = 16'hcd91;
mem_array[9394] = 16'h3e88;
mem_array[9397] = 16'heb46;
mem_array[9396] = 16'hbe34;
mem_array[9399] = 16'ha994;
mem_array[9398] = 16'hbdaa;
mem_array[9401] = 16'h7aa5;
mem_array[9400] = 16'h3ec8;
mem_array[9403] = 16'h2451;
mem_array[9402] = 16'h3e31;
mem_array[9405] = 16'h4b52;
mem_array[9404] = 16'hbf0e;
mem_array[9407] = 16'hcd65;
mem_array[9406] = 16'h3d5f;
mem_array[9409] = 16'h470a;
mem_array[9408] = 16'hbe2b;
mem_array[9411] = 16'hc0f5;
mem_array[9410] = 16'hbf28;
mem_array[9413] = 16'h7494;
mem_array[9412] = 16'h3e0b;
mem_array[9415] = 16'h0247;
mem_array[9414] = 16'hbe37;
mem_array[9417] = 16'h7f68;
mem_array[9416] = 16'h3e2d;
mem_array[9419] = 16'h3f16;
mem_array[9418] = 16'hbead;
mem_array[9421] = 16'h206b;
mem_array[9420] = 16'hbdfc;
mem_array[9423] = 16'h23f0;
mem_array[9422] = 16'hbf8c;
mem_array[9425] = 16'hd185;
mem_array[9424] = 16'hbe2d;
mem_array[9427] = 16'h6952;
mem_array[9426] = 16'h3d17;
mem_array[9429] = 16'hd526;
mem_array[9428] = 16'hbf26;
mem_array[9431] = 16'ha623;
mem_array[9430] = 16'h3e26;
mem_array[9433] = 16'hb52c;
mem_array[9432] = 16'hbe06;
mem_array[9435] = 16'h1e7a;
mem_array[9434] = 16'hbe49;
mem_array[9437] = 16'h28a2;
mem_array[9436] = 16'hbe29;
mem_array[9439] = 16'hab90;
mem_array[9438] = 16'hbda2;
mem_array[9441] = 16'h6421;
mem_array[9440] = 16'h3ba0;
mem_array[9443] = 16'h5e60;
mem_array[9442] = 16'h3b61;
mem_array[9445] = 16'h5c43;
mem_array[9444] = 16'h3d8c;
mem_array[9447] = 16'h8f10;
mem_array[9446] = 16'h3d52;
mem_array[9449] = 16'h1f3b;
mem_array[9448] = 16'h3e0c;
mem_array[9451] = 16'h7c91;
mem_array[9450] = 16'hbe28;
mem_array[9453] = 16'h6ffa;
mem_array[9452] = 16'hbe83;
mem_array[9455] = 16'h7596;
mem_array[9454] = 16'h3ec9;
mem_array[9457] = 16'hfe88;
mem_array[9456] = 16'hbf23;
mem_array[9459] = 16'hb7a5;
mem_array[9458] = 16'h3e7c;
mem_array[9461] = 16'hc390;
mem_array[9460] = 16'h3ead;
mem_array[9463] = 16'h844b;
mem_array[9462] = 16'h3e7c;
mem_array[9465] = 16'hb59b;
mem_array[9464] = 16'hbd78;
mem_array[9467] = 16'h7689;
mem_array[9466] = 16'hbc84;
mem_array[9469] = 16'hfcce;
mem_array[9468] = 16'hbd9d;
mem_array[9471] = 16'h5cec;
mem_array[9470] = 16'hbf14;
mem_array[9473] = 16'h748b;
mem_array[9472] = 16'h3e7b;
mem_array[9475] = 16'he77a;
mem_array[9474] = 16'hbe62;
mem_array[9477] = 16'hb9eb;
mem_array[9476] = 16'hbdc2;
mem_array[9479] = 16'h7ad6;
mem_array[9478] = 16'hbd87;
mem_array[9481] = 16'h5804;
mem_array[9480] = 16'h3c77;
mem_array[9483] = 16'h123b;
mem_array[9482] = 16'hbfc7;
mem_array[9485] = 16'h023b;
mem_array[9484] = 16'hbe46;
mem_array[9487] = 16'h2c44;
mem_array[9486] = 16'h3c23;
mem_array[9489] = 16'h2c3a;
mem_array[9488] = 16'hbebb;
mem_array[9491] = 16'h7ef4;
mem_array[9490] = 16'h3d98;
mem_array[9493] = 16'hc8e4;
mem_array[9492] = 16'hbc6b;
mem_array[9495] = 16'hf0cc;
mem_array[9494] = 16'h3e17;
mem_array[9497] = 16'h886d;
mem_array[9496] = 16'h3e13;
mem_array[9499] = 16'h03f3;
mem_array[9498] = 16'hbed7;
mem_array[9501] = 16'hf73b;
mem_array[9500] = 16'hbd3d;
mem_array[9503] = 16'h8bfb;
mem_array[9502] = 16'hbce1;
mem_array[9505] = 16'h052f;
mem_array[9504] = 16'hbdc1;
mem_array[9507] = 16'ha4f3;
mem_array[9506] = 16'h3d08;
mem_array[9509] = 16'h7345;
mem_array[9508] = 16'h3e39;
mem_array[9511] = 16'h6588;
mem_array[9510] = 16'hbd52;
mem_array[9513] = 16'hdbbc;
mem_array[9512] = 16'h3e82;
mem_array[9515] = 16'h896f;
mem_array[9514] = 16'h3e08;
mem_array[9517] = 16'hd740;
mem_array[9516] = 16'hbe8e;
mem_array[9519] = 16'h863e;
mem_array[9518] = 16'h3e9f;
mem_array[9521] = 16'h044a;
mem_array[9520] = 16'hbf06;
mem_array[9523] = 16'hc71a;
mem_array[9522] = 16'hbe6f;
mem_array[9525] = 16'hf5df;
mem_array[9524] = 16'hbbc9;
mem_array[9527] = 16'h6a6d;
mem_array[9526] = 16'hbdf0;
mem_array[9529] = 16'h22ce;
mem_array[9528] = 16'hbdf1;
mem_array[9531] = 16'h9160;
mem_array[9530] = 16'hbf4c;
mem_array[9533] = 16'hc0a9;
mem_array[9532] = 16'h3e6a;
mem_array[9535] = 16'h4c4e;
mem_array[9534] = 16'hbf01;
mem_array[9537] = 16'h6110;
mem_array[9536] = 16'h3d9c;
mem_array[9539] = 16'h896e;
mem_array[9538] = 16'h3e2a;
mem_array[9541] = 16'h8de9;
mem_array[9540] = 16'h3e24;
mem_array[9543] = 16'h4243;
mem_array[9542] = 16'hbf90;
mem_array[9545] = 16'h48e0;
mem_array[9544] = 16'hbe3c;
mem_array[9547] = 16'hb2b4;
mem_array[9546] = 16'h3e9a;
mem_array[9549] = 16'hf239;
mem_array[9548] = 16'hbdbf;
mem_array[9551] = 16'hdf0d;
mem_array[9550] = 16'h3e38;
mem_array[9553] = 16'h0d6f;
mem_array[9552] = 16'hbcb6;
mem_array[9555] = 16'h68af;
mem_array[9554] = 16'h3e3b;
mem_array[9557] = 16'h7286;
mem_array[9556] = 16'h3edf;
mem_array[9559] = 16'hb0dd;
mem_array[9558] = 16'hbec4;
mem_array[9561] = 16'hdef3;
mem_array[9560] = 16'hbd6c;
mem_array[9563] = 16'h14e4;
mem_array[9562] = 16'h3d85;
mem_array[9565] = 16'h0876;
mem_array[9564] = 16'h3b9c;
mem_array[9567] = 16'he282;
mem_array[9566] = 16'h3ea0;
mem_array[9569] = 16'h72eb;
mem_array[9568] = 16'h3e89;
mem_array[9571] = 16'h5b20;
mem_array[9570] = 16'hbe3d;
mem_array[9573] = 16'h3fbd;
mem_array[9572] = 16'h3d1f;
mem_array[9575] = 16'h655b;
mem_array[9574] = 16'h3e33;
mem_array[9577] = 16'hd031;
mem_array[9576] = 16'hbd60;
mem_array[9579] = 16'h7ac3;
mem_array[9578] = 16'h3ed3;
mem_array[9581] = 16'hcc51;
mem_array[9580] = 16'hbea1;
mem_array[9583] = 16'h77e3;
mem_array[9582] = 16'hbea9;
mem_array[9585] = 16'h735d;
mem_array[9584] = 16'h3c3f;
mem_array[9587] = 16'hb5ac;
mem_array[9586] = 16'hbd04;
mem_array[9589] = 16'h036a;
mem_array[9588] = 16'hbeb1;
mem_array[9591] = 16'he605;
mem_array[9590] = 16'hbfed;
mem_array[9593] = 16'h8f47;
mem_array[9592] = 16'h3e4a;
mem_array[9595] = 16'hcce5;
mem_array[9594] = 16'hbf2e;
mem_array[9597] = 16'h9e38;
mem_array[9596] = 16'h3edb;
mem_array[9599] = 16'hc90d;
mem_array[9598] = 16'h3e76;
mem_array[9601] = 16'h931e;
mem_array[9600] = 16'hbcab;
mem_array[9603] = 16'h4681;
mem_array[9602] = 16'hbf7b;
mem_array[9605] = 16'h744a;
mem_array[9604] = 16'hbe6c;
mem_array[9607] = 16'hf371;
mem_array[9606] = 16'h3bbf;
mem_array[9609] = 16'h8fee;
mem_array[9608] = 16'hbda8;
mem_array[9611] = 16'hd173;
mem_array[9610] = 16'h3e11;
mem_array[9613] = 16'h8fda;
mem_array[9612] = 16'h3cee;
mem_array[9615] = 16'hfe8a;
mem_array[9614] = 16'hbdd8;
mem_array[9617] = 16'h8e39;
mem_array[9616] = 16'h3eac;
mem_array[9619] = 16'hc407;
mem_array[9618] = 16'hbfd9;
mem_array[9621] = 16'h5cae;
mem_array[9620] = 16'hbd4f;
mem_array[9623] = 16'ha028;
mem_array[9622] = 16'hbdd7;
mem_array[9625] = 16'hd6b9;
mem_array[9624] = 16'hbdae;
mem_array[9627] = 16'h9b59;
mem_array[9626] = 16'h3e3e;
mem_array[9629] = 16'hc0c4;
mem_array[9628] = 16'h3e9e;
mem_array[9631] = 16'h2192;
mem_array[9630] = 16'hbe4a;
mem_array[9633] = 16'hc788;
mem_array[9632] = 16'h3ec2;
mem_array[9635] = 16'h00fa;
mem_array[9634] = 16'h3e73;
mem_array[9637] = 16'h7eb8;
mem_array[9636] = 16'hbef5;
mem_array[9639] = 16'h5d4a;
mem_array[9638] = 16'hbb9a;
mem_array[9641] = 16'h5c37;
mem_array[9640] = 16'hbe45;
mem_array[9643] = 16'h1214;
mem_array[9642] = 16'hbd3b;
mem_array[9645] = 16'h60a9;
mem_array[9644] = 16'h3f12;
mem_array[9647] = 16'h92c1;
mem_array[9646] = 16'hbdba;
mem_array[9649] = 16'h1ae1;
mem_array[9648] = 16'h3cc0;
mem_array[9651] = 16'hef9a;
mem_array[9650] = 16'hbf63;
mem_array[9653] = 16'hbdb6;
mem_array[9652] = 16'h3ecf;
mem_array[9655] = 16'h2df2;
mem_array[9654] = 16'hbee1;
mem_array[9657] = 16'h3247;
mem_array[9656] = 16'hbe35;
mem_array[9659] = 16'h1a25;
mem_array[9658] = 16'hbe95;
mem_array[9661] = 16'hbf5f;
mem_array[9660] = 16'h3e22;
mem_array[9663] = 16'h8516;
mem_array[9662] = 16'hbe8a;
mem_array[9665] = 16'hb2a7;
mem_array[9664] = 16'hbe88;
mem_array[9667] = 16'h0074;
mem_array[9666] = 16'hbc5e;
mem_array[9669] = 16'h31a5;
mem_array[9668] = 16'hbb04;
mem_array[9671] = 16'h27f6;
mem_array[9670] = 16'h3e26;
mem_array[9673] = 16'h060e;
mem_array[9672] = 16'hbea4;
mem_array[9675] = 16'h4e82;
mem_array[9674] = 16'hbd92;
mem_array[9677] = 16'h12b2;
mem_array[9676] = 16'hbefc;
mem_array[9679] = 16'h1147;
mem_array[9678] = 16'hbfb6;
mem_array[9681] = 16'h6e49;
mem_array[9680] = 16'h3d1f;
mem_array[9683] = 16'he050;
mem_array[9682] = 16'hbdcc;
mem_array[9685] = 16'hc6ef;
mem_array[9684] = 16'hbe8b;
mem_array[9687] = 16'h4c59;
mem_array[9686] = 16'h3eb6;
mem_array[9689] = 16'h3d33;
mem_array[9688] = 16'hbd5f;
mem_array[9691] = 16'hf4a5;
mem_array[9690] = 16'hbd59;
mem_array[9693] = 16'h649e;
mem_array[9692] = 16'h3e65;
mem_array[9695] = 16'h91b4;
mem_array[9694] = 16'h3ea2;
mem_array[9697] = 16'hc54f;
mem_array[9696] = 16'hbed4;
mem_array[9699] = 16'hfe7b;
mem_array[9698] = 16'h3e42;
mem_array[9701] = 16'h8bf7;
mem_array[9700] = 16'h3e22;
mem_array[9703] = 16'hcaae;
mem_array[9702] = 16'hbcae;
mem_array[9705] = 16'h4310;
mem_array[9704] = 16'h3d8d;
mem_array[9707] = 16'hc4cc;
mem_array[9706] = 16'hbdd6;
mem_array[9709] = 16'h8e4f;
mem_array[9708] = 16'hbf13;
mem_array[9711] = 16'h59e3;
mem_array[9710] = 16'hbf7d;
mem_array[9713] = 16'hae80;
mem_array[9712] = 16'h3ef9;
mem_array[9715] = 16'ha469;
mem_array[9714] = 16'hbe90;
mem_array[9717] = 16'ha2e0;
mem_array[9716] = 16'h3e82;
mem_array[9719] = 16'h8709;
mem_array[9718] = 16'hbd00;
mem_array[9721] = 16'h3bf6;
mem_array[9720] = 16'h3f41;
mem_array[9723] = 16'h52ed;
mem_array[9722] = 16'hbf3c;
mem_array[9725] = 16'h240c;
mem_array[9724] = 16'h3d5a;
mem_array[9727] = 16'h96a4;
mem_array[9726] = 16'h3e18;
mem_array[9729] = 16'hca56;
mem_array[9728] = 16'hbce3;
mem_array[9731] = 16'h546b;
mem_array[9730] = 16'h3ec0;
mem_array[9733] = 16'h604f;
mem_array[9732] = 16'hbf1d;
mem_array[9735] = 16'hc279;
mem_array[9734] = 16'hbbe4;
mem_array[9737] = 16'ha6f7;
mem_array[9736] = 16'hbf67;
mem_array[9739] = 16'h6a29;
mem_array[9738] = 16'hbe82;
mem_array[9741] = 16'h29a5;
mem_array[9740] = 16'h3dad;
mem_array[9743] = 16'h6e33;
mem_array[9742] = 16'h3cfb;
mem_array[9745] = 16'hfff9;
mem_array[9744] = 16'hbec2;
mem_array[9747] = 16'h9c42;
mem_array[9746] = 16'h3e9b;
mem_array[9749] = 16'hbba3;
mem_array[9748] = 16'h3ee1;
mem_array[9751] = 16'h3ba5;
mem_array[9750] = 16'hbdb2;
mem_array[9753] = 16'hb73d;
mem_array[9752] = 16'h3c4e;
mem_array[9755] = 16'he441;
mem_array[9754] = 16'hbc62;
mem_array[9757] = 16'h7b2f;
mem_array[9756] = 16'hbf56;
mem_array[9759] = 16'h760e;
mem_array[9758] = 16'h3ed3;
mem_array[9761] = 16'heac5;
mem_array[9760] = 16'h3d96;
mem_array[9763] = 16'hbc2e;
mem_array[9762] = 16'hbdbd;
mem_array[9765] = 16'h2ef4;
mem_array[9764] = 16'hbe56;
mem_array[9767] = 16'h2d9e;
mem_array[9766] = 16'hbdf0;
mem_array[9769] = 16'h5c2c;
mem_array[9768] = 16'hbe98;
mem_array[9771] = 16'hfee2;
mem_array[9770] = 16'h3e33;
mem_array[9773] = 16'hf5e0;
mem_array[9772] = 16'h3f08;
mem_array[9775] = 16'h3bd3;
mem_array[9774] = 16'hbc76;
mem_array[9777] = 16'hc3bb;
mem_array[9776] = 16'h3e1c;
mem_array[9779] = 16'h5bf2;
mem_array[9778] = 16'h3c08;
mem_array[9781] = 16'h1d74;
mem_array[9780] = 16'h3e80;
mem_array[9783] = 16'hb6a5;
mem_array[9782] = 16'hbdb1;
mem_array[9785] = 16'hf432;
mem_array[9784] = 16'h3f12;
mem_array[9787] = 16'h3895;
mem_array[9786] = 16'h3da3;
mem_array[9789] = 16'h731d;
mem_array[9788] = 16'hbe59;
mem_array[9791] = 16'he664;
mem_array[9790] = 16'h3f20;
mem_array[9793] = 16'h1bde;
mem_array[9792] = 16'hbf25;
mem_array[9795] = 16'hbc0b;
mem_array[9794] = 16'hbe7c;
mem_array[9797] = 16'h6896;
mem_array[9796] = 16'hbfc1;
mem_array[9799] = 16'h0bc8;
mem_array[9798] = 16'hbec6;
mem_array[9801] = 16'h363e;
mem_array[9800] = 16'h3d80;
mem_array[9803] = 16'hf828;
mem_array[9802] = 16'h3d87;
mem_array[9805] = 16'h3a9e;
mem_array[9804] = 16'hbedf;
mem_array[9807] = 16'h1820;
mem_array[9806] = 16'h3d12;
mem_array[9809] = 16'h47ed;
mem_array[9808] = 16'h3e2a;
mem_array[9811] = 16'hc7ca;
mem_array[9810] = 16'hbe65;
mem_array[9813] = 16'hd136;
mem_array[9812] = 16'hbd7f;
mem_array[9815] = 16'h4e96;
mem_array[9814] = 16'hbe03;
mem_array[9817] = 16'hb655;
mem_array[9816] = 16'hbe65;
mem_array[9819] = 16'h2826;
mem_array[9818] = 16'h3f33;
mem_array[9821] = 16'h2bd4;
mem_array[9820] = 16'h3ec8;
mem_array[9823] = 16'h1265;
mem_array[9822] = 16'hbe9d;
mem_array[9825] = 16'h92b5;
mem_array[9824] = 16'hbe91;
mem_array[9827] = 16'h9d1c;
mem_array[9826] = 16'hbeab;
mem_array[9829] = 16'h8e37;
mem_array[9828] = 16'hbe62;
mem_array[9831] = 16'h13ed;
mem_array[9830] = 16'hbeda;
mem_array[9833] = 16'h02d3;
mem_array[9832] = 16'h3eb3;
mem_array[9835] = 16'hbeb8;
mem_array[9834] = 16'h3de7;
mem_array[9837] = 16'ha57a;
mem_array[9836] = 16'hbf23;
mem_array[9839] = 16'h3787;
mem_array[9838] = 16'h3ef3;
mem_array[9841] = 16'h96fa;
mem_array[9840] = 16'h3e02;
mem_array[9843] = 16'hf9c9;
mem_array[9842] = 16'h3e70;
mem_array[9845] = 16'h4d7e;
mem_array[9844] = 16'hbed1;
mem_array[9847] = 16'h3cfb;
mem_array[9846] = 16'hbeb4;
mem_array[9849] = 16'h9e40;
mem_array[9848] = 16'h3e1e;
mem_array[9851] = 16'h2f69;
mem_array[9850] = 16'h3ee8;
mem_array[9853] = 16'h3d77;
mem_array[9852] = 16'hbf25;
mem_array[9855] = 16'h4ef4;
mem_array[9854] = 16'hbf04;
mem_array[9857] = 16'hd631;
mem_array[9856] = 16'hbf24;
mem_array[9859] = 16'h5192;
mem_array[9858] = 16'h3e0c;
mem_array[9861] = 16'h49bf;
mem_array[9860] = 16'hbd80;
mem_array[9863] = 16'hf01d;
mem_array[9862] = 16'hbb48;
mem_array[9865] = 16'h1553;
mem_array[9864] = 16'h3b67;
mem_array[9867] = 16'hd9d7;
mem_array[9866] = 16'hbf75;
mem_array[9869] = 16'h9678;
mem_array[9868] = 16'hbed1;
mem_array[9871] = 16'h261b;
mem_array[9870] = 16'hbe80;
mem_array[9873] = 16'h5fc8;
mem_array[9872] = 16'h3d53;
mem_array[9875] = 16'hb06e;
mem_array[9874] = 16'hbe82;
mem_array[9877] = 16'h5673;
mem_array[9876] = 16'hbe07;
mem_array[9879] = 16'hb66b;
mem_array[9878] = 16'h3e11;
mem_array[9881] = 16'h4e9e;
mem_array[9880] = 16'h3ea1;
mem_array[9883] = 16'h96ad;
mem_array[9882] = 16'hbe68;
mem_array[9885] = 16'h262c;
mem_array[9884] = 16'hbebb;
mem_array[9887] = 16'h2a41;
mem_array[9886] = 16'hbe78;
mem_array[9889] = 16'haf8e;
mem_array[9888] = 16'hbf96;
mem_array[9891] = 16'h6ae6;
mem_array[9890] = 16'hbe45;
mem_array[9893] = 16'h170e;
mem_array[9892] = 16'h3d0f;
mem_array[9895] = 16'h9990;
mem_array[9894] = 16'hbdbc;
mem_array[9897] = 16'h6b4c;
mem_array[9896] = 16'hbf3b;
mem_array[9899] = 16'hc792;
mem_array[9898] = 16'h3ed5;
mem_array[9901] = 16'hb615;
mem_array[9900] = 16'hbee5;
mem_array[9903] = 16'h21c3;
mem_array[9902] = 16'h3f51;
mem_array[9905] = 16'h0aa4;
mem_array[9904] = 16'hbde1;
mem_array[9907] = 16'h604b;
mem_array[9906] = 16'hbfcc;
mem_array[9909] = 16'h8c35;
mem_array[9908] = 16'hbe44;
mem_array[9911] = 16'h76ee;
mem_array[9910] = 16'h3da6;
mem_array[9913] = 16'h6e9e;
mem_array[9912] = 16'h3e23;
mem_array[9915] = 16'h090c;
mem_array[9914] = 16'hbee6;
mem_array[9917] = 16'h86de;
mem_array[9916] = 16'h3f1f;
mem_array[9919] = 16'h7c76;
mem_array[9918] = 16'hbd77;
mem_array[9921] = 16'h41c5;
mem_array[9920] = 16'hbd8e;
mem_array[9923] = 16'hf8ab;
mem_array[9922] = 16'h3d52;
mem_array[9925] = 16'hc17d;
mem_array[9924] = 16'hbf35;
mem_array[9927] = 16'h747d;
mem_array[9926] = 16'h3f65;
mem_array[9929] = 16'h5d03;
mem_array[9928] = 16'hbf01;
mem_array[9931] = 16'hb877;
mem_array[9930] = 16'hbd2d;
mem_array[9933] = 16'h283f;
mem_array[9932] = 16'hbec1;
mem_array[9935] = 16'hbdc2;
mem_array[9934] = 16'hbdd0;
mem_array[9937] = 16'h5829;
mem_array[9936] = 16'h3eb6;
mem_array[9939] = 16'h29d3;
mem_array[9938] = 16'h3f7f;
mem_array[9941] = 16'ha560;
mem_array[9940] = 16'h3e71;
mem_array[9943] = 16'h67ee;
mem_array[9942] = 16'hbe18;
mem_array[9945] = 16'h2014;
mem_array[9944] = 16'hbf43;
mem_array[9947] = 16'h26f1;
mem_array[9946] = 16'hbef6;
mem_array[9949] = 16'he970;
mem_array[9948] = 16'hbf72;
mem_array[9951] = 16'h9d01;
mem_array[9950] = 16'hbea5;
mem_array[9953] = 16'h2e85;
mem_array[9952] = 16'hbe46;
mem_array[9955] = 16'h15d0;
mem_array[9954] = 16'h3f25;
mem_array[9957] = 16'hf703;
mem_array[9956] = 16'h3edc;
mem_array[9959] = 16'h03da;
mem_array[9958] = 16'hbf0c;
mem_array[9961] = 16'h088b;
mem_array[9960] = 16'hbe47;
mem_array[9963] = 16'hca84;
mem_array[9962] = 16'h3f16;
mem_array[9965] = 16'h79a3;
mem_array[9964] = 16'hbf06;
mem_array[9967] = 16'ha139;
mem_array[9966] = 16'hbfbb;
mem_array[9969] = 16'hcdde;
mem_array[9968] = 16'h3e90;
mem_array[9971] = 16'h7f62;
mem_array[9970] = 16'h3f20;
mem_array[9973] = 16'he1bd;
mem_array[9972] = 16'h3d59;
mem_array[9975] = 16'h90a6;
mem_array[9974] = 16'h3f1a;
mem_array[9977] = 16'he4fc;
mem_array[9976] = 16'hbd43;
mem_array[9979] = 16'hbf8d;
mem_array[9978] = 16'hbd2d;
mem_array[9981] = 16'hd824;
mem_array[9980] = 16'hbc1e;
mem_array[9983] = 16'h6de9;
mem_array[9982] = 16'hbd67;
mem_array[9985] = 16'h944b;
mem_array[9984] = 16'h3e95;
mem_array[9987] = 16'h6601;
mem_array[9986] = 16'hbde1;
mem_array[9989] = 16'h193e;
mem_array[9988] = 16'hbda9;
mem_array[9991] = 16'hbb0f;
mem_array[9990] = 16'hbf58;
mem_array[9993] = 16'h1796;
mem_array[9992] = 16'hbf1d;
mem_array[9995] = 16'h249b;
mem_array[9994] = 16'hbed7;
mem_array[9997] = 16'hd054;
mem_array[9996] = 16'h3f11;
mem_array[9999] = 16'hd102;
mem_array[9998] = 16'h3eb7;
mem_array[10001] = 16'ha447;
mem_array[10000] = 16'hbfbf;
mem_array[10003] = 16'h9796;
mem_array[10002] = 16'h3ee6;
mem_array[10005] = 16'h3f06;
mem_array[10004] = 16'hbf20;
mem_array[10007] = 16'h0061;
mem_array[10006] = 16'h3c52;
mem_array[10009] = 16'h4613;
mem_array[10008] = 16'hbd92;
mem_array[10011] = 16'h4e30;
mem_array[10010] = 16'hbe5b;
mem_array[10013] = 16'h05bb;
mem_array[10012] = 16'h3f3a;
mem_array[10015] = 16'hb187;
mem_array[10014] = 16'h3f5e;
mem_array[10017] = 16'h5486;
mem_array[10016] = 16'hbd9b;
mem_array[10019] = 16'hdc0f;
mem_array[10018] = 16'hbf2b;
mem_array[10021] = 16'hffbe;
mem_array[10020] = 16'hbdc8;
mem_array[10023] = 16'h3920;
mem_array[10022] = 16'h3ea5;
mem_array[10025] = 16'heece;
mem_array[10024] = 16'hbe54;
mem_array[10027] = 16'hebd7;
mem_array[10026] = 16'hbf41;
mem_array[10029] = 16'he682;
mem_array[10028] = 16'hbb09;
mem_array[10031] = 16'he5ea;
mem_array[10030] = 16'h3e2e;
mem_array[10033] = 16'h914c;
mem_array[10032] = 16'h3de0;
mem_array[10035] = 16'h63c3;
mem_array[10034] = 16'h3e88;
mem_array[10037] = 16'hf021;
mem_array[10036] = 16'h3c15;
mem_array[10039] = 16'h1277;
mem_array[10038] = 16'h3cf2;
mem_array[10041] = 16'h3aed;
mem_array[10040] = 16'hbca2;
mem_array[10043] = 16'h70b1;
mem_array[10042] = 16'h3c7d;
mem_array[10045] = 16'hb752;
mem_array[10044] = 16'h3f45;
mem_array[10047] = 16'h166b;
mem_array[10046] = 16'hbe49;
mem_array[10049] = 16'h5156;
mem_array[10048] = 16'hbda0;
mem_array[10051] = 16'hf90c;
mem_array[10050] = 16'hbf2a;
mem_array[10053] = 16'h33e0;
mem_array[10052] = 16'hbf06;
mem_array[10055] = 16'hf6bf;
mem_array[10054] = 16'hbc18;
mem_array[10057] = 16'ha167;
mem_array[10056] = 16'hbe50;
mem_array[10059] = 16'h14b9;
mem_array[10058] = 16'h3cad;
mem_array[10061] = 16'h0977;
mem_array[10060] = 16'h3e3a;
mem_array[10063] = 16'he35d;
mem_array[10062] = 16'h3db3;
mem_array[10065] = 16'he509;
mem_array[10064] = 16'h3e0e;
mem_array[10067] = 16'hb609;
mem_array[10066] = 16'h3f30;
mem_array[10069] = 16'h4f78;
mem_array[10068] = 16'hbe36;
mem_array[10071] = 16'h794d;
mem_array[10070] = 16'hbcd7;
mem_array[10073] = 16'hff8f;
mem_array[10072] = 16'hbecb;
mem_array[10075] = 16'hf810;
mem_array[10074] = 16'h3eac;
mem_array[10077] = 16'he8ab;
mem_array[10076] = 16'h3d5f;
mem_array[10079] = 16'h660e;
mem_array[10078] = 16'h3ebd;
mem_array[10081] = 16'hccac;
mem_array[10080] = 16'hbcbc;
mem_array[10083] = 16'h2182;
mem_array[10082] = 16'hbdc7;
mem_array[10085] = 16'hcd0a;
mem_array[10084] = 16'hbd65;
mem_array[10087] = 16'h9c65;
mem_array[10086] = 16'hbdbd;
mem_array[10089] = 16'hd6c7;
mem_array[10088] = 16'h3d23;
mem_array[10091] = 16'h58b3;
mem_array[10090] = 16'h3c84;
mem_array[10093] = 16'hf500;
mem_array[10092] = 16'hbd92;
mem_array[10095] = 16'h2e09;
mem_array[10094] = 16'hbd96;
mem_array[10097] = 16'h2fe6;
mem_array[10096] = 16'h3dc0;
mem_array[10099] = 16'h7d24;
mem_array[10098] = 16'hbc94;
mem_array[10101] = 16'h2aa0;
mem_array[10100] = 16'h3d86;
mem_array[10103] = 16'h2c6c;
mem_array[10102] = 16'hbcda;
mem_array[10105] = 16'h3243;
mem_array[10104] = 16'hbc5d;
mem_array[10107] = 16'h55e7;
mem_array[10106] = 16'hbb47;
mem_array[10109] = 16'ha1d1;
mem_array[10108] = 16'h3dd7;
mem_array[10111] = 16'h51fa;
mem_array[10110] = 16'hbb23;
mem_array[10113] = 16'h689e;
mem_array[10112] = 16'hbb61;
mem_array[10115] = 16'h4ce2;
mem_array[10114] = 16'hbc84;
mem_array[10117] = 16'h4b72;
mem_array[10116] = 16'h3c88;
mem_array[10119] = 16'h50dd;
mem_array[10118] = 16'hbd93;
mem_array[10121] = 16'h798c;
mem_array[10120] = 16'h3d30;
mem_array[10123] = 16'h182c;
mem_array[10122] = 16'hbb9c;
mem_array[10125] = 16'h79db;
mem_array[10124] = 16'hbd1e;
mem_array[10127] = 16'hf812;
mem_array[10126] = 16'h3d12;
mem_array[10129] = 16'h7643;
mem_array[10128] = 16'h3cbf;
mem_array[10131] = 16'hc3dd;
mem_array[10130] = 16'h3da6;
mem_array[10133] = 16'h1a4c;
mem_array[10132] = 16'hbd5f;
mem_array[10135] = 16'hd362;
mem_array[10134] = 16'hbd4f;
mem_array[10137] = 16'h554a;
mem_array[10136] = 16'h3c36;
mem_array[10139] = 16'hd509;
mem_array[10138] = 16'hbb6d;
mem_array[10141] = 16'h3749;
mem_array[10140] = 16'h3c81;
mem_array[10143] = 16'hf324;
mem_array[10142] = 16'h3c0c;
mem_array[10145] = 16'heb7e;
mem_array[10144] = 16'h3d28;
mem_array[10147] = 16'h4434;
mem_array[10146] = 16'h3de0;
mem_array[10149] = 16'hb116;
mem_array[10148] = 16'hbc94;
mem_array[10151] = 16'h34d7;
mem_array[10150] = 16'hbae5;
mem_array[10153] = 16'hb9f3;
mem_array[10152] = 16'h3d92;
mem_array[10155] = 16'ha988;
mem_array[10154] = 16'h3dd1;
mem_array[10157] = 16'hde23;
mem_array[10156] = 16'h3d06;
mem_array[10159] = 16'hd1ca;
mem_array[10158] = 16'h3d31;
mem_array[10161] = 16'h4c0b;
mem_array[10160] = 16'h3d26;
mem_array[10163] = 16'hd2eb;
mem_array[10162] = 16'hbdc5;
mem_array[10165] = 16'h44c8;
mem_array[10164] = 16'h3d6c;
mem_array[10167] = 16'h8c2a;
mem_array[10166] = 16'h3c24;
mem_array[10169] = 16'h929d;
mem_array[10168] = 16'hbbc0;
mem_array[10171] = 16'h77ab;
mem_array[10170] = 16'h3ca9;
mem_array[10173] = 16'hd844;
mem_array[10172] = 16'h3c79;
mem_array[10175] = 16'h6bdf;
mem_array[10174] = 16'h3d9c;
mem_array[10177] = 16'h9eff;
mem_array[10176] = 16'h3cf8;
mem_array[10179] = 16'h5dc0;
mem_array[10178] = 16'h3bf8;
mem_array[10181] = 16'h8ca1;
mem_array[10180] = 16'hbe34;
mem_array[10183] = 16'h7cb2;
mem_array[10182] = 16'h3e29;
mem_array[10185] = 16'h40e4;
mem_array[10184] = 16'h3b49;
mem_array[10187] = 16'h0111;
mem_array[10186] = 16'hbf20;
mem_array[10189] = 16'hef39;
mem_array[10188] = 16'h3f15;
mem_array[10191] = 16'h51b0;
mem_array[10190] = 16'hbd02;
mem_array[10193] = 16'h1835;
mem_array[10192] = 16'h3ef0;
mem_array[10195] = 16'h84ef;
mem_array[10194] = 16'h3d0e;
mem_array[10197] = 16'ha0a6;
mem_array[10196] = 16'h3d47;
mem_array[10199] = 16'h5a72;
mem_array[10198] = 16'hbc8e;
mem_array[10201] = 16'h53f6;
mem_array[10200] = 16'hbdbc;
mem_array[10203] = 16'h5aa5;
mem_array[10202] = 16'h3d9c;
mem_array[10205] = 16'h88d0;
mem_array[10204] = 16'h3bdd;
mem_array[10207] = 16'h7e8f;
mem_array[10206] = 16'hbef8;
mem_array[10209] = 16'h08d2;
mem_array[10208] = 16'h3dcf;
mem_array[10211] = 16'h4eb9;
mem_array[10210] = 16'h3f10;
mem_array[10213] = 16'h2aea;
mem_array[10212] = 16'h3f9b;
mem_array[10215] = 16'he29b;
mem_array[10214] = 16'h3e7e;
mem_array[10217] = 16'h82ff;
mem_array[10216] = 16'h3c03;
mem_array[10219] = 16'h4bdc;
mem_array[10218] = 16'h3ec0;
mem_array[10221] = 16'h31da;
mem_array[10220] = 16'h3d1f;
mem_array[10223] = 16'hbb31;
mem_array[10222] = 16'h3c88;
mem_array[10225] = 16'h4f5e;
mem_array[10224] = 16'hbf0c;
mem_array[10227] = 16'h53da;
mem_array[10226] = 16'h3e56;
mem_array[10229] = 16'h2f00;
mem_array[10228] = 16'h3f09;
mem_array[10231] = 16'h9c7e;
mem_array[10230] = 16'hbebe;
mem_array[10233] = 16'hca5b;
mem_array[10232] = 16'h3e43;
mem_array[10235] = 16'h3834;
mem_array[10234] = 16'hbe1d;
mem_array[10237] = 16'h803e;
mem_array[10236] = 16'h3eb6;
mem_array[10239] = 16'h8878;
mem_array[10238] = 16'h3ece;
mem_array[10241] = 16'hbb64;
mem_array[10240] = 16'h3bdb;
mem_array[10243] = 16'he4fb;
mem_array[10242] = 16'hbda1;
mem_array[10245] = 16'h7163;
mem_array[10244] = 16'hbda0;
mem_array[10247] = 16'h2445;
mem_array[10246] = 16'hbed4;
mem_array[10249] = 16'h9679;
mem_array[10248] = 16'h3f26;
mem_array[10251] = 16'h2cf3;
mem_array[10250] = 16'h3eb8;
mem_array[10253] = 16'h2112;
mem_array[10252] = 16'h3e09;
mem_array[10255] = 16'hab5c;
mem_array[10254] = 16'h3e98;
mem_array[10257] = 16'h1b32;
mem_array[10256] = 16'h3efc;
mem_array[10259] = 16'hbf10;
mem_array[10258] = 16'hbdd0;
mem_array[10261] = 16'h02e7;
mem_array[10260] = 16'h3f08;
mem_array[10263] = 16'hb9f9;
mem_array[10262] = 16'h3f20;
mem_array[10265] = 16'h7d5d;
mem_array[10264] = 16'hbf57;
mem_array[10267] = 16'h10a3;
mem_array[10266] = 16'hbf73;
mem_array[10269] = 16'h6df6;
mem_array[10268] = 16'h3ed4;
mem_array[10271] = 16'ha7cd;
mem_array[10270] = 16'h3e6d;
mem_array[10273] = 16'haeed;
mem_array[10272] = 16'h3f1d;
mem_array[10275] = 16'h51e4;
mem_array[10274] = 16'h3ee0;
mem_array[10277] = 16'haf63;
mem_array[10276] = 16'hbeb2;
mem_array[10279] = 16'hfca7;
mem_array[10278] = 16'hbe47;
mem_array[10281] = 16'h67a9;
mem_array[10280] = 16'h3dba;
mem_array[10283] = 16'hbc4b;
mem_array[10282] = 16'h3d55;
mem_array[10285] = 16'h20a3;
mem_array[10284] = 16'hbe55;
mem_array[10287] = 16'h69ee;
mem_array[10286] = 16'hbf16;
mem_array[10289] = 16'h4f10;
mem_array[10288] = 16'hbf40;
mem_array[10291] = 16'h72b3;
mem_array[10290] = 16'h3e08;
mem_array[10293] = 16'h027c;
mem_array[10292] = 16'h3eaf;
mem_array[10295] = 16'hf183;
mem_array[10294] = 16'h3e55;
mem_array[10297] = 16'h3c8f;
mem_array[10296] = 16'h3fad;
mem_array[10299] = 16'h5d92;
mem_array[10298] = 16'h3f17;
mem_array[10301] = 16'h297e;
mem_array[10300] = 16'hbe6f;
mem_array[10303] = 16'h78b6;
mem_array[10302] = 16'h3ed7;
mem_array[10305] = 16'h0a84;
mem_array[10304] = 16'hbe1c;
mem_array[10307] = 16'h68cc;
mem_array[10306] = 16'hbdb1;
mem_array[10309] = 16'h3986;
mem_array[10308] = 16'h3ddc;
mem_array[10311] = 16'h5576;
mem_array[10310] = 16'h3fad;
mem_array[10313] = 16'h7fdf;
mem_array[10312] = 16'h3ea3;
mem_array[10315] = 16'h0150;
mem_array[10314] = 16'h3eeb;
mem_array[10317] = 16'h39d1;
mem_array[10316] = 16'h3ec4;
mem_array[10319] = 16'h9b73;
mem_array[10318] = 16'hbeab;
mem_array[10321] = 16'h45cc;
mem_array[10320] = 16'h3f0b;
mem_array[10323] = 16'h2f89;
mem_array[10322] = 16'h3f19;
mem_array[10325] = 16'h6c0a;
mem_array[10324] = 16'h3d1c;
mem_array[10327] = 16'h4847;
mem_array[10326] = 16'h3ebd;
mem_array[10329] = 16'hfa24;
mem_array[10328] = 16'h3ebc;
mem_array[10331] = 16'h8bb4;
mem_array[10330] = 16'hbed4;
mem_array[10333] = 16'hb969;
mem_array[10332] = 16'h3ecb;
mem_array[10335] = 16'h6f7a;
mem_array[10334] = 16'h3f65;
mem_array[10337] = 16'hfad2;
mem_array[10336] = 16'h3ee3;
mem_array[10339] = 16'ha0e5;
mem_array[10338] = 16'hbd37;
mem_array[10341] = 16'h7eaf;
mem_array[10340] = 16'h3cb1;
mem_array[10343] = 16'h2f86;
mem_array[10342] = 16'h3cb8;
mem_array[10345] = 16'h31e0;
mem_array[10344] = 16'hbf38;
mem_array[10347] = 16'h39e4;
mem_array[10346] = 16'h3f02;
mem_array[10349] = 16'h418a;
mem_array[10348] = 16'hbe62;
mem_array[10351] = 16'hf44f;
mem_array[10350] = 16'hbf56;
mem_array[10353] = 16'hf7d5;
mem_array[10352] = 16'h3f29;
mem_array[10355] = 16'he43b;
mem_array[10354] = 16'hbefc;
mem_array[10357] = 16'h7bce;
mem_array[10356] = 16'hbefa;
mem_array[10359] = 16'h0e02;
mem_array[10358] = 16'h3e2e;
mem_array[10361] = 16'h27b0;
mem_array[10360] = 16'h3e1b;
mem_array[10363] = 16'h514b;
mem_array[10362] = 16'h3e96;
mem_array[10365] = 16'hab32;
mem_array[10364] = 16'hbe1a;
mem_array[10367] = 16'h140e;
mem_array[10366] = 16'h3d7b;
mem_array[10369] = 16'h07db;
mem_array[10368] = 16'hbe83;
mem_array[10371] = 16'h526a;
mem_array[10370] = 16'h3f21;
mem_array[10373] = 16'h6c22;
mem_array[10372] = 16'h3e3d;
mem_array[10375] = 16'hf4b0;
mem_array[10374] = 16'h3db6;
mem_array[10377] = 16'h345e;
mem_array[10376] = 16'h3df5;
mem_array[10379] = 16'h543e;
mem_array[10378] = 16'h3d52;
mem_array[10381] = 16'h2b09;
mem_array[10380] = 16'h3b96;
mem_array[10383] = 16'haa1b;
mem_array[10382] = 16'h3f14;
mem_array[10385] = 16'h6701;
mem_array[10384] = 16'hbe65;
mem_array[10387] = 16'hca6c;
mem_array[10386] = 16'h3e11;
mem_array[10389] = 16'h7092;
mem_array[10388] = 16'hbd77;
mem_array[10391] = 16'he938;
mem_array[10390] = 16'hbf96;
mem_array[10393] = 16'hd699;
mem_array[10392] = 16'h3f0d;
mem_array[10395] = 16'h8e71;
mem_array[10394] = 16'hbe17;
mem_array[10397] = 16'h8f3c;
mem_array[10396] = 16'hbde7;
mem_array[10399] = 16'h7c6f;
mem_array[10398] = 16'hbf2c;
mem_array[10401] = 16'hb79b;
mem_array[10400] = 16'h3db4;
mem_array[10403] = 16'hbf65;
mem_array[10402] = 16'hbbd7;
mem_array[10405] = 16'hc36a;
mem_array[10404] = 16'hbeb8;
mem_array[10407] = 16'h6625;
mem_array[10406] = 16'h3e10;
mem_array[10409] = 16'h6cb5;
mem_array[10408] = 16'hbe54;
mem_array[10411] = 16'h0738;
mem_array[10410] = 16'hbe8e;
mem_array[10413] = 16'h8481;
mem_array[10412] = 16'hbec3;
mem_array[10415] = 16'hfd5e;
mem_array[10414] = 16'h3e94;
mem_array[10417] = 16'hd601;
mem_array[10416] = 16'hbe44;
mem_array[10419] = 16'haf3c;
mem_array[10418] = 16'h3ec9;
mem_array[10421] = 16'h9f46;
mem_array[10420] = 16'h3f45;
mem_array[10423] = 16'h870b;
mem_array[10422] = 16'h3e69;
mem_array[10425] = 16'h8d09;
mem_array[10424] = 16'hbf80;
mem_array[10427] = 16'h075a;
mem_array[10426] = 16'hbd44;
mem_array[10429] = 16'ha015;
mem_array[10428] = 16'hbe84;
mem_array[10431] = 16'hb564;
mem_array[10430] = 16'h3f78;
mem_array[10433] = 16'h23c6;
mem_array[10432] = 16'hbed4;
mem_array[10435] = 16'h1a94;
mem_array[10434] = 16'hbcc8;
mem_array[10437] = 16'h08b5;
mem_array[10436] = 16'hbdbe;
mem_array[10439] = 16'h84b8;
mem_array[10438] = 16'h3ee0;
mem_array[10441] = 16'hf621;
mem_array[10440] = 16'hbf15;
mem_array[10443] = 16'hef0e;
mem_array[10442] = 16'hbe11;
mem_array[10445] = 16'hf59b;
mem_array[10444] = 16'h3d82;
mem_array[10447] = 16'hf4d7;
mem_array[10446] = 16'hbdab;
mem_array[10449] = 16'hd75f;
mem_array[10448] = 16'h3e28;
mem_array[10451] = 16'h2b80;
mem_array[10450] = 16'hbe42;
mem_array[10453] = 16'h939b;
mem_array[10452] = 16'h3ead;
mem_array[10455] = 16'h4cfe;
mem_array[10454] = 16'hbec2;
mem_array[10457] = 16'hfab0;
mem_array[10456] = 16'h3e33;
mem_array[10459] = 16'hbc0d;
mem_array[10458] = 16'hbebb;
mem_array[10461] = 16'haa2a;
mem_array[10460] = 16'hbb30;
mem_array[10463] = 16'hd184;
mem_array[10462] = 16'h3c98;
mem_array[10465] = 16'h5333;
mem_array[10464] = 16'h3cbf;
mem_array[10467] = 16'h9a9b;
mem_array[10466] = 16'h3df5;
mem_array[10469] = 16'hef3b;
mem_array[10468] = 16'hbeb9;
mem_array[10471] = 16'hadfd;
mem_array[10470] = 16'hbd82;
mem_array[10473] = 16'h0b3b;
mem_array[10472] = 16'hbcf2;
mem_array[10475] = 16'h6174;
mem_array[10474] = 16'h3e0f;
mem_array[10477] = 16'hc1ba;
mem_array[10476] = 16'h3e6e;
mem_array[10479] = 16'haf09;
mem_array[10478] = 16'h3c5a;
mem_array[10481] = 16'hb5ac;
mem_array[10480] = 16'hbd5f;
mem_array[10483] = 16'ha467;
mem_array[10482] = 16'h3e6f;
mem_array[10485] = 16'h1aab;
mem_array[10484] = 16'hbf93;
mem_array[10487] = 16'h1926;
mem_array[10486] = 16'hbe8e;
mem_array[10489] = 16'h85b7;
mem_array[10488] = 16'hbdf3;
mem_array[10491] = 16'hebc9;
mem_array[10490] = 16'h3eab;
mem_array[10493] = 16'haaf5;
mem_array[10492] = 16'hbef4;
mem_array[10495] = 16'hefbe;
mem_array[10494] = 16'hbecc;
mem_array[10497] = 16'h9f9a;
mem_array[10496] = 16'h3edf;
mem_array[10499] = 16'h04f5;
mem_array[10498] = 16'h3d37;
mem_array[10501] = 16'hb506;
mem_array[10500] = 16'h3d68;
mem_array[10503] = 16'hc310;
mem_array[10502] = 16'h3c25;
mem_array[10505] = 16'h3d6a;
mem_array[10504] = 16'h3d06;
mem_array[10507] = 16'h0dd2;
mem_array[10506] = 16'h3db8;
mem_array[10509] = 16'h1bbe;
mem_array[10508] = 16'h3ee6;
mem_array[10511] = 16'h03e3;
mem_array[10510] = 16'hbf37;
mem_array[10513] = 16'h03d8;
mem_array[10512] = 16'h3ead;
mem_array[10515] = 16'h7dae;
mem_array[10514] = 16'hbcdd;
mem_array[10517] = 16'h18b2;
mem_array[10516] = 16'h3e84;
mem_array[10519] = 16'h404c;
mem_array[10518] = 16'hbf58;
mem_array[10521] = 16'hd43c;
mem_array[10520] = 16'hbc84;
mem_array[10523] = 16'hfa7f;
mem_array[10522] = 16'h3c4d;
mem_array[10525] = 16'h260a;
mem_array[10524] = 16'h3d0a;
mem_array[10527] = 16'hcd8f;
mem_array[10526] = 16'hbe0d;
mem_array[10529] = 16'h00f1;
mem_array[10528] = 16'hbf04;
mem_array[10531] = 16'h63af;
mem_array[10530] = 16'hbe32;
mem_array[10533] = 16'hfd2a;
mem_array[10532] = 16'h3cee;
mem_array[10535] = 16'h9722;
mem_array[10534] = 16'h3c78;
mem_array[10537] = 16'hf715;
mem_array[10536] = 16'h3ebc;
mem_array[10539] = 16'hfacf;
mem_array[10538] = 16'hbd9b;
mem_array[10541] = 16'hd47c;
mem_array[10540] = 16'h3c2f;
mem_array[10543] = 16'h1542;
mem_array[10542] = 16'hbd73;
mem_array[10545] = 16'hcd77;
mem_array[10544] = 16'hbf00;
mem_array[10547] = 16'h2748;
mem_array[10546] = 16'h3e8b;
mem_array[10549] = 16'h776a;
mem_array[10548] = 16'h3d0a;
mem_array[10551] = 16'h897b;
mem_array[10550] = 16'h3e69;
mem_array[10553] = 16'h6769;
mem_array[10552] = 16'hbd23;
mem_array[10555] = 16'h0898;
mem_array[10554] = 16'hbf1b;
mem_array[10557] = 16'ha8f5;
mem_array[10556] = 16'h3e2d;
mem_array[10559] = 16'h2e05;
mem_array[10558] = 16'h3d16;
mem_array[10561] = 16'hbf89;
mem_array[10560] = 16'hbec2;
mem_array[10563] = 16'hf815;
mem_array[10562] = 16'h3a0f;
mem_array[10565] = 16'h4b58;
mem_array[10564] = 16'h3e33;
mem_array[10567] = 16'hd3aa;
mem_array[10566] = 16'hbe33;
mem_array[10569] = 16'h4710;
mem_array[10568] = 16'h3ed3;
mem_array[10571] = 16'h11d1;
mem_array[10570] = 16'hbeb9;
mem_array[10573] = 16'h8817;
mem_array[10572] = 16'h3e50;
mem_array[10575] = 16'h7601;
mem_array[10574] = 16'h3e35;
mem_array[10577] = 16'h53e5;
mem_array[10576] = 16'hbd5a;
mem_array[10579] = 16'h4c25;
mem_array[10578] = 16'hbebc;
mem_array[10581] = 16'h4267;
mem_array[10580] = 16'h3db6;
mem_array[10583] = 16'hf006;
mem_array[10582] = 16'hbcfc;
mem_array[10585] = 16'h1ed0;
mem_array[10584] = 16'h3de2;
mem_array[10587] = 16'hb6da;
mem_array[10586] = 16'h3d28;
mem_array[10589] = 16'ha700;
mem_array[10588] = 16'hbdcd;
mem_array[10591] = 16'h5276;
mem_array[10590] = 16'hbd53;
mem_array[10593] = 16'h02dd;
mem_array[10592] = 16'h3e89;
mem_array[10595] = 16'hd1de;
mem_array[10594] = 16'h3d93;
mem_array[10597] = 16'hd18f;
mem_array[10596] = 16'hbcd1;
mem_array[10599] = 16'hcc02;
mem_array[10598] = 16'h3e69;
mem_array[10601] = 16'h2f6a;
mem_array[10600] = 16'hbe94;
mem_array[10603] = 16'h0cf3;
mem_array[10602] = 16'h3e85;
mem_array[10605] = 16'h9fe5;
mem_array[10604] = 16'h3da3;
mem_array[10607] = 16'h8f09;
mem_array[10606] = 16'hbd7e;
mem_array[10609] = 16'hd8ef;
mem_array[10608] = 16'hbe2e;
mem_array[10611] = 16'h29e7;
mem_array[10610] = 16'h3e80;
mem_array[10613] = 16'h801f;
mem_array[10612] = 16'h3eab;
mem_array[10615] = 16'hc9f4;
mem_array[10614] = 16'hbf3e;
mem_array[10617] = 16'h992d;
mem_array[10616] = 16'hbea2;
mem_array[10619] = 16'h6c97;
mem_array[10618] = 16'hbeb5;
mem_array[10621] = 16'h7139;
mem_array[10620] = 16'h3ed7;
mem_array[10623] = 16'h2df1;
mem_array[10622] = 16'hbf50;
mem_array[10625] = 16'h6e57;
mem_array[10624] = 16'h3eae;
mem_array[10627] = 16'h2ed2;
mem_array[10626] = 16'hbf06;
mem_array[10629] = 16'h07ba;
mem_array[10628] = 16'h3db3;
mem_array[10631] = 16'he523;
mem_array[10630] = 16'hbedb;
mem_array[10633] = 16'hc261;
mem_array[10632] = 16'h3e86;
mem_array[10635] = 16'hd27a;
mem_array[10634] = 16'hbda5;
mem_array[10637] = 16'hed05;
mem_array[10636] = 16'h3d2a;
mem_array[10639] = 16'h5b97;
mem_array[10638] = 16'hbeed;
mem_array[10641] = 16'hfdce;
mem_array[10640] = 16'hbdca;
mem_array[10643] = 16'h04ea;
mem_array[10642] = 16'hbca3;
mem_array[10645] = 16'hbcec;
mem_array[10644] = 16'hbe5b;
mem_array[10647] = 16'hb930;
mem_array[10646] = 16'h3d43;
mem_array[10649] = 16'h0915;
mem_array[10648] = 16'hbd2b;
mem_array[10651] = 16'h3463;
mem_array[10650] = 16'hbdbe;
mem_array[10653] = 16'hc87a;
mem_array[10652] = 16'h3dfd;
mem_array[10655] = 16'hec46;
mem_array[10654] = 16'h3ebf;
mem_array[10657] = 16'h310c;
mem_array[10656] = 16'h3dda;
mem_array[10659] = 16'h429a;
mem_array[10658] = 16'h3e41;
mem_array[10661] = 16'h5834;
mem_array[10660] = 16'h3e66;
mem_array[10663] = 16'h2c9d;
mem_array[10662] = 16'hbd41;
mem_array[10665] = 16'h7851;
mem_array[10664] = 16'h3ea2;
mem_array[10667] = 16'h6811;
mem_array[10666] = 16'hbe67;
mem_array[10669] = 16'h6bbc;
mem_array[10668] = 16'h3e84;
mem_array[10671] = 16'h5feb;
mem_array[10670] = 16'h3edd;
mem_array[10673] = 16'hedbf;
mem_array[10672] = 16'hbd79;
mem_array[10675] = 16'h8827;
mem_array[10674] = 16'hbec3;
mem_array[10677] = 16'hdfd5;
mem_array[10676] = 16'hbdda;
mem_array[10679] = 16'h4a0b;
mem_array[10678] = 16'hbe67;
mem_array[10681] = 16'h9ce9;
mem_array[10680] = 16'h3e8a;
mem_array[10683] = 16'h3916;
mem_array[10682] = 16'hbf1d;
mem_array[10685] = 16'h4f02;
mem_array[10684] = 16'h3d79;
mem_array[10687] = 16'h92ca;
mem_array[10686] = 16'hbdab;
mem_array[10689] = 16'h14e1;
mem_array[10688] = 16'h3dac;
mem_array[10691] = 16'h1d87;
mem_array[10690] = 16'h3d25;
mem_array[10693] = 16'h4fc4;
mem_array[10692] = 16'h3d17;
mem_array[10695] = 16'h5f51;
mem_array[10694] = 16'h3ea1;
mem_array[10697] = 16'h3622;
mem_array[10696] = 16'h3e00;
mem_array[10699] = 16'h745f;
mem_array[10698] = 16'hbf69;
mem_array[10701] = 16'h6c60;
mem_array[10700] = 16'hbc9a;
mem_array[10703] = 16'hc16f;
mem_array[10702] = 16'h3d4a;
mem_array[10705] = 16'hc50f;
mem_array[10704] = 16'hbdea;
mem_array[10707] = 16'h28fa;
mem_array[10706] = 16'hbe05;
mem_array[10709] = 16'h8055;
mem_array[10708] = 16'hbe2d;
mem_array[10711] = 16'h612f;
mem_array[10710] = 16'h3e53;
mem_array[10713] = 16'hcd60;
mem_array[10712] = 16'hbdff;
mem_array[10715] = 16'h6f20;
mem_array[10714] = 16'hbe95;
mem_array[10717] = 16'hb2b6;
mem_array[10716] = 16'hbe44;
mem_array[10719] = 16'h282a;
mem_array[10718] = 16'hbd61;
mem_array[10721] = 16'h4338;
mem_array[10720] = 16'hbedb;
mem_array[10723] = 16'h44ad;
mem_array[10722] = 16'h3eae;
mem_array[10725] = 16'hbbf7;
mem_array[10724] = 16'h3e14;
mem_array[10727] = 16'h0e00;
mem_array[10726] = 16'h3d31;
mem_array[10729] = 16'h450a;
mem_array[10728] = 16'h3e0d;
mem_array[10731] = 16'h262f;
mem_array[10730] = 16'hbdcf;
mem_array[10733] = 16'haba5;
mem_array[10732] = 16'h3e66;
mem_array[10735] = 16'h2c67;
mem_array[10734] = 16'hbe08;
mem_array[10737] = 16'h6448;
mem_array[10736] = 16'hbe21;
mem_array[10739] = 16'h6626;
mem_array[10738] = 16'hbf2c;
mem_array[10741] = 16'h1798;
mem_array[10740] = 16'h3e6f;
mem_array[10743] = 16'hc135;
mem_array[10742] = 16'h3d0d;
mem_array[10745] = 16'hbc7b;
mem_array[10744] = 16'h3d70;
mem_array[10747] = 16'h0ae5;
mem_array[10746] = 16'h3c9c;
mem_array[10749] = 16'h55c7;
mem_array[10748] = 16'h3ecd;
mem_array[10751] = 16'h1ac5;
mem_array[10750] = 16'h3e85;
mem_array[10753] = 16'h74d0;
mem_array[10752] = 16'h3e15;
mem_array[10755] = 16'he969;
mem_array[10754] = 16'h3da2;
mem_array[10757] = 16'hd105;
mem_array[10756] = 16'h3ef4;
mem_array[10759] = 16'h69a5;
mem_array[10758] = 16'hbe56;
mem_array[10761] = 16'h10ea;
mem_array[10760] = 16'hbd22;
mem_array[10763] = 16'h76bb;
mem_array[10762] = 16'hbd2d;
mem_array[10765] = 16'hc501;
mem_array[10764] = 16'h3ca2;
mem_array[10767] = 16'h640e;
mem_array[10766] = 16'h3e34;
mem_array[10769] = 16'h1b7b;
mem_array[10768] = 16'hbbdb;
mem_array[10771] = 16'h43e2;
mem_array[10770] = 16'h3e68;
mem_array[10773] = 16'h425b;
mem_array[10772] = 16'hbea6;
mem_array[10775] = 16'h3dc1;
mem_array[10774] = 16'hbe43;
mem_array[10777] = 16'h0ce0;
mem_array[10776] = 16'h3da3;
mem_array[10779] = 16'h1724;
mem_array[10778] = 16'hbdd4;
mem_array[10781] = 16'hc7f3;
mem_array[10780] = 16'hbf2c;
mem_array[10783] = 16'hb7bf;
mem_array[10782] = 16'h3cb0;
mem_array[10785] = 16'hbde4;
mem_array[10784] = 16'hbe36;
mem_array[10787] = 16'he0e9;
mem_array[10786] = 16'hbdee;
mem_array[10789] = 16'hfc42;
mem_array[10788] = 16'h3cd7;
mem_array[10791] = 16'hf268;
mem_array[10790] = 16'h3e37;
mem_array[10793] = 16'h674b;
mem_array[10792] = 16'hbc32;
mem_array[10795] = 16'hecf4;
mem_array[10794] = 16'hbe23;
mem_array[10797] = 16'h7023;
mem_array[10796] = 16'hbe2f;
mem_array[10799] = 16'hfec6;
mem_array[10798] = 16'hbf24;
mem_array[10801] = 16'hc8a2;
mem_array[10800] = 16'hbf6d;
mem_array[10803] = 16'h9226;
mem_array[10802] = 16'h3db7;
mem_array[10805] = 16'hffd3;
mem_array[10804] = 16'h3df2;
mem_array[10807] = 16'h2500;
mem_array[10806] = 16'h3c7d;
mem_array[10809] = 16'h4065;
mem_array[10808] = 16'h3eb0;
mem_array[10811] = 16'h0695;
mem_array[10810] = 16'hbdd6;
mem_array[10813] = 16'h25ee;
mem_array[10812] = 16'h3ddc;
mem_array[10815] = 16'hbad5;
mem_array[10814] = 16'h3e85;
mem_array[10817] = 16'hcf51;
mem_array[10816] = 16'h3e6d;
mem_array[10819] = 16'h554a;
mem_array[10818] = 16'hbc96;
mem_array[10821] = 16'hc1c9;
mem_array[10820] = 16'hbca4;
mem_array[10823] = 16'he8f7;
mem_array[10822] = 16'hbd48;
mem_array[10825] = 16'h3105;
mem_array[10824] = 16'hbcbb;
mem_array[10827] = 16'hd120;
mem_array[10826] = 16'h3b04;
mem_array[10829] = 16'h529c;
mem_array[10828] = 16'hbd96;
mem_array[10831] = 16'h969e;
mem_array[10830] = 16'hbe0c;
mem_array[10833] = 16'h7d5a;
mem_array[10832] = 16'hbd6a;
mem_array[10835] = 16'ha5ef;
mem_array[10834] = 16'hbeb6;
mem_array[10837] = 16'hd2dd;
mem_array[10836] = 16'hbb96;
mem_array[10839] = 16'hdfb6;
mem_array[10838] = 16'hbeb3;
mem_array[10841] = 16'hfd5b;
mem_array[10840] = 16'hbe65;
mem_array[10843] = 16'h597f;
mem_array[10842] = 16'h3d04;
mem_array[10845] = 16'h8e83;
mem_array[10844] = 16'hbca7;
mem_array[10847] = 16'h0c5f;
mem_array[10846] = 16'hbe31;
mem_array[10849] = 16'h1d76;
mem_array[10848] = 16'hbe44;
mem_array[10851] = 16'hd18c;
mem_array[10850] = 16'h3ecd;
mem_array[10853] = 16'h611b;
mem_array[10852] = 16'h3cfe;
mem_array[10855] = 16'he66b;
mem_array[10854] = 16'h3e36;
mem_array[10857] = 16'hf012;
mem_array[10856] = 16'h3e0f;
mem_array[10859] = 16'he26d;
mem_array[10858] = 16'hbec5;
mem_array[10861] = 16'he1a2;
mem_array[10860] = 16'hbf95;
mem_array[10863] = 16'h8234;
mem_array[10862] = 16'hbe09;
mem_array[10865] = 16'h58d2;
mem_array[10864] = 16'h3d15;
mem_array[10867] = 16'h316d;
mem_array[10866] = 16'h3db7;
mem_array[10869] = 16'hf984;
mem_array[10868] = 16'h3d01;
mem_array[10871] = 16'h0058;
mem_array[10870] = 16'hbe3d;
mem_array[10873] = 16'hc147;
mem_array[10872] = 16'h3e71;
mem_array[10875] = 16'h9591;
mem_array[10874] = 16'h3e4e;
mem_array[10877] = 16'h050d;
mem_array[10876] = 16'h3e18;
mem_array[10879] = 16'h3b2e;
mem_array[10878] = 16'hbe25;
mem_array[10881] = 16'hd18e;
mem_array[10880] = 16'hbaab;
mem_array[10883] = 16'h7f24;
mem_array[10882] = 16'hbd23;
mem_array[10885] = 16'h800e;
mem_array[10884] = 16'h3d83;
mem_array[10887] = 16'h23aa;
mem_array[10886] = 16'h3e29;
mem_array[10889] = 16'h210d;
mem_array[10888] = 16'hbdd1;
mem_array[10891] = 16'h3698;
mem_array[10890] = 16'hbe02;
mem_array[10893] = 16'hcb61;
mem_array[10892] = 16'hbda6;
mem_array[10895] = 16'ha29c;
mem_array[10894] = 16'hbed2;
mem_array[10897] = 16'hec48;
mem_array[10896] = 16'hbd04;
mem_array[10899] = 16'hdfce;
mem_array[10898] = 16'hbe2f;
mem_array[10901] = 16'he49f;
mem_array[10900] = 16'hbe63;
mem_array[10903] = 16'headb;
mem_array[10902] = 16'hbca1;
mem_array[10905] = 16'hd8e9;
mem_array[10904] = 16'hbf13;
mem_array[10907] = 16'h24ec;
mem_array[10906] = 16'h3c49;
mem_array[10909] = 16'h283e;
mem_array[10908] = 16'hbd8e;
mem_array[10911] = 16'h6eec;
mem_array[10910] = 16'hbe82;
mem_array[10913] = 16'h7cfe;
mem_array[10912] = 16'hbbb8;
mem_array[10915] = 16'h4421;
mem_array[10914] = 16'h3e62;
mem_array[10917] = 16'hb3c5;
mem_array[10916] = 16'h3d00;
mem_array[10919] = 16'ha2e2;
mem_array[10918] = 16'hbea4;
mem_array[10921] = 16'hdd66;
mem_array[10920] = 16'hbea2;
mem_array[10923] = 16'h31eb;
mem_array[10922] = 16'hbe23;
mem_array[10925] = 16'h2673;
mem_array[10924] = 16'h3d29;
mem_array[10927] = 16'h22bd;
mem_array[10926] = 16'h3e86;
mem_array[10929] = 16'h6ab7;
mem_array[10928] = 16'h3cf6;
mem_array[10931] = 16'h58fb;
mem_array[10930] = 16'hbd9f;
mem_array[10933] = 16'h5c8e;
mem_array[10932] = 16'h3e4e;
mem_array[10935] = 16'h8946;
mem_array[10934] = 16'h3c4c;
mem_array[10937] = 16'ha5e5;
mem_array[10936] = 16'h3d08;
mem_array[10939] = 16'ha5f0;
mem_array[10938] = 16'hbdd4;
mem_array[10941] = 16'h5b18;
mem_array[10940] = 16'hbd96;
mem_array[10943] = 16'h0f42;
mem_array[10942] = 16'hbd5f;
mem_array[10945] = 16'hb23d;
mem_array[10944] = 16'hbe86;
mem_array[10947] = 16'h00f1;
mem_array[10946] = 16'h3e0d;
mem_array[10949] = 16'h9410;
mem_array[10948] = 16'hbe37;
mem_array[10951] = 16'h4905;
mem_array[10950] = 16'hbdea;
mem_array[10953] = 16'hd245;
mem_array[10952] = 16'hbe14;
mem_array[10955] = 16'h6c07;
mem_array[10954] = 16'hbf2e;
mem_array[10957] = 16'h7e4e;
mem_array[10956] = 16'h3dc8;
mem_array[10959] = 16'h35a4;
mem_array[10958] = 16'h3e35;
mem_array[10961] = 16'hc640;
mem_array[10960] = 16'hbe09;
mem_array[10963] = 16'h4953;
mem_array[10962] = 16'h3c85;
mem_array[10965] = 16'h3019;
mem_array[10964] = 16'hbd5a;
mem_array[10967] = 16'habd5;
mem_array[10966] = 16'hbe81;
mem_array[10969] = 16'h84af;
mem_array[10968] = 16'hbd97;
mem_array[10971] = 16'h1cb3;
mem_array[10970] = 16'hbf0e;
mem_array[10973] = 16'h3848;
mem_array[10972] = 16'h3d6e;
mem_array[10975] = 16'h8876;
mem_array[10974] = 16'h3da0;
mem_array[10977] = 16'h8d38;
mem_array[10976] = 16'hbdfb;
mem_array[10979] = 16'hbb29;
mem_array[10978] = 16'hbf12;
mem_array[10981] = 16'hde67;
mem_array[10980] = 16'hbed2;
mem_array[10983] = 16'h7dc3;
mem_array[10982] = 16'hbe4b;
mem_array[10985] = 16'h3247;
mem_array[10984] = 16'h3cb3;
mem_array[10987] = 16'h9900;
mem_array[10986] = 16'hbc41;
mem_array[10989] = 16'h4605;
mem_array[10988] = 16'hbe45;
mem_array[10991] = 16'ha335;
mem_array[10990] = 16'hbe95;
mem_array[10993] = 16'hf2cd;
mem_array[10992] = 16'hbcf5;
mem_array[10995] = 16'hf352;
mem_array[10994] = 16'h3c95;
mem_array[10997] = 16'h07a5;
mem_array[10996] = 16'hbe7c;
mem_array[10999] = 16'hf715;
mem_array[10998] = 16'h3d55;
mem_array[11001] = 16'hcf7f;
mem_array[11000] = 16'hbc96;
mem_array[11003] = 16'h4e0f;
mem_array[11002] = 16'h3bab;
mem_array[11005] = 16'h4189;
mem_array[11004] = 16'hbe99;
mem_array[11007] = 16'h4b77;
mem_array[11006] = 16'h3e42;
mem_array[11009] = 16'h8131;
mem_array[11008] = 16'hbda7;
mem_array[11011] = 16'hb15a;
mem_array[11010] = 16'hbd9b;
mem_array[11013] = 16'h21af;
mem_array[11012] = 16'hbe8a;
mem_array[11015] = 16'h4dee;
mem_array[11014] = 16'hbfde;
mem_array[11017] = 16'h8bd7;
mem_array[11016] = 16'hbd0d;
mem_array[11019] = 16'hca7d;
mem_array[11018] = 16'hbee8;
mem_array[11021] = 16'h6471;
mem_array[11020] = 16'hbe59;
mem_array[11023] = 16'hf812;
mem_array[11022] = 16'hbdd0;
mem_array[11025] = 16'heeeb;
mem_array[11024] = 16'hbe5e;
mem_array[11027] = 16'h008c;
mem_array[11026] = 16'hbd9b;
mem_array[11029] = 16'h5392;
mem_array[11028] = 16'h3d45;
mem_array[11031] = 16'h209f;
mem_array[11030] = 16'hbe23;
mem_array[11033] = 16'h58df;
mem_array[11032] = 16'h3e5e;
mem_array[11035] = 16'h9f7f;
mem_array[11034] = 16'hbe92;
mem_array[11037] = 16'h6b12;
mem_array[11036] = 16'h3e11;
mem_array[11039] = 16'h22ab;
mem_array[11038] = 16'hbef8;
mem_array[11041] = 16'hb3f6;
mem_array[11040] = 16'hbe28;
mem_array[11043] = 16'ha0da;
mem_array[11042] = 16'hbeb4;
mem_array[11045] = 16'ha5da;
mem_array[11044] = 16'h3e3d;
mem_array[11047] = 16'h7db3;
mem_array[11046] = 16'hbe36;
mem_array[11049] = 16'h8681;
mem_array[11048] = 16'hbe48;
mem_array[11051] = 16'h0cf8;
mem_array[11050] = 16'hbe06;
mem_array[11053] = 16'h4224;
mem_array[11052] = 16'hbe93;
mem_array[11055] = 16'h129d;
mem_array[11054] = 16'h3e9b;
mem_array[11057] = 16'he854;
mem_array[11056] = 16'hbdbe;
mem_array[11059] = 16'h6932;
mem_array[11058] = 16'hbe86;
mem_array[11061] = 16'h1e7e;
mem_array[11060] = 16'hbd5d;
mem_array[11063] = 16'h5646;
mem_array[11062] = 16'hbd9b;
mem_array[11065] = 16'h5772;
mem_array[11064] = 16'hbeae;
mem_array[11067] = 16'h3568;
mem_array[11066] = 16'h3e0c;
mem_array[11069] = 16'h834b;
mem_array[11068] = 16'h3cae;
mem_array[11071] = 16'h9b11;
mem_array[11070] = 16'hbd9a;
mem_array[11073] = 16'h03a7;
mem_array[11072] = 16'hbd87;
mem_array[11075] = 16'h7184;
mem_array[11074] = 16'hbe6f;
mem_array[11077] = 16'hf92e;
mem_array[11076] = 16'hbd76;
mem_array[11079] = 16'h3293;
mem_array[11078] = 16'hbec3;
mem_array[11081] = 16'hd7a1;
mem_array[11080] = 16'h3d21;
mem_array[11083] = 16'hcab8;
mem_array[11082] = 16'h3e11;
mem_array[11085] = 16'hb6c2;
mem_array[11084] = 16'hbf1d;
mem_array[11087] = 16'he9e1;
mem_array[11086] = 16'h3d17;
mem_array[11089] = 16'h92e9;
mem_array[11088] = 16'h3e10;
mem_array[11091] = 16'h4abd;
mem_array[11090] = 16'hbd01;
mem_array[11093] = 16'h3ee4;
mem_array[11092] = 16'h3e5c;
mem_array[11095] = 16'h05ed;
mem_array[11094] = 16'hbea9;
mem_array[11097] = 16'h6002;
mem_array[11096] = 16'h3e54;
mem_array[11099] = 16'h411a;
mem_array[11098] = 16'hbee9;
mem_array[11101] = 16'hd26e;
mem_array[11100] = 16'hbe1b;
mem_array[11103] = 16'h30f6;
mem_array[11102] = 16'h3e7c;
mem_array[11105] = 16'h4eb6;
mem_array[11104] = 16'h3d6c;
mem_array[11107] = 16'he0de;
mem_array[11106] = 16'hbd47;
mem_array[11109] = 16'ha318;
mem_array[11108] = 16'hba54;
mem_array[11111] = 16'h17fb;
mem_array[11110] = 16'h3e4c;
mem_array[11113] = 16'hbd42;
mem_array[11112] = 16'hbd98;
mem_array[11115] = 16'hba59;
mem_array[11114] = 16'h3c9b;
mem_array[11117] = 16'h5904;
mem_array[11116] = 16'h3ebd;
mem_array[11119] = 16'h83e4;
mem_array[11118] = 16'hbed6;
mem_array[11121] = 16'h7f09;
mem_array[11120] = 16'h3bb9;
mem_array[11123] = 16'h50e6;
mem_array[11122] = 16'hbda2;
mem_array[11125] = 16'h7dd1;
mem_array[11124] = 16'hbf0e;
mem_array[11127] = 16'haa84;
mem_array[11126] = 16'h3d3e;
mem_array[11129] = 16'h24a2;
mem_array[11128] = 16'h3db4;
mem_array[11131] = 16'h7a89;
mem_array[11130] = 16'hbcb8;
mem_array[11133] = 16'h483b;
mem_array[11132] = 16'h3df2;
mem_array[11135] = 16'hc598;
mem_array[11134] = 16'h3d86;
mem_array[11137] = 16'h10ff;
mem_array[11136] = 16'h3f0f;
mem_array[11139] = 16'hbd18;
mem_array[11138] = 16'hbeb0;
mem_array[11141] = 16'h22ea;
mem_array[11140] = 16'hbe19;
mem_array[11143] = 16'h2df5;
mem_array[11142] = 16'h3e40;
mem_array[11145] = 16'h6e03;
mem_array[11144] = 16'hbe28;
mem_array[11147] = 16'he616;
mem_array[11146] = 16'hbea9;
mem_array[11149] = 16'ha7ed;
mem_array[11148] = 16'hbdc1;
mem_array[11151] = 16'h6cab;
mem_array[11150] = 16'hbd45;
mem_array[11153] = 16'hb1f1;
mem_array[11152] = 16'h3e05;
mem_array[11155] = 16'h98cf;
mem_array[11154] = 16'hbdc6;
mem_array[11157] = 16'h2764;
mem_array[11156] = 16'h3da8;
mem_array[11159] = 16'hd9e9;
mem_array[11158] = 16'hbee9;
mem_array[11161] = 16'h29fc;
mem_array[11160] = 16'hbe03;
mem_array[11163] = 16'h28cc;
mem_array[11162] = 16'h3ecc;
mem_array[11165] = 16'h4e16;
mem_array[11164] = 16'hbe08;
mem_array[11167] = 16'hfbc9;
mem_array[11166] = 16'h3e08;
mem_array[11169] = 16'hbeec;
mem_array[11168] = 16'h3cfd;
mem_array[11171] = 16'h56d3;
mem_array[11170] = 16'h3e72;
mem_array[11173] = 16'hf36e;
mem_array[11172] = 16'h3d05;
mem_array[11175] = 16'hfe72;
mem_array[11174] = 16'h3cad;
mem_array[11177] = 16'h70b4;
mem_array[11176] = 16'h3e16;
mem_array[11179] = 16'h301f;
mem_array[11178] = 16'hbdd8;
mem_array[11181] = 16'h2838;
mem_array[11180] = 16'hbdb0;
mem_array[11183] = 16'hfbe2;
mem_array[11182] = 16'hbd0d;
mem_array[11185] = 16'h94fc;
mem_array[11184] = 16'hbe99;
mem_array[11187] = 16'h70a7;
mem_array[11186] = 16'h3e6a;
mem_array[11189] = 16'had18;
mem_array[11188] = 16'h3db6;
mem_array[11191] = 16'h0065;
mem_array[11190] = 16'hbd22;
mem_array[11193] = 16'hfc05;
mem_array[11192] = 16'h3ede;
mem_array[11195] = 16'hb526;
mem_array[11194] = 16'h3dbc;
mem_array[11197] = 16'hfa88;
mem_array[11196] = 16'h3eac;
mem_array[11199] = 16'h33f7;
mem_array[11198] = 16'hbef8;
mem_array[11201] = 16'h9e72;
mem_array[11200] = 16'hbeff;
mem_array[11203] = 16'h35c1;
mem_array[11202] = 16'h3c13;
mem_array[11205] = 16'h7423;
mem_array[11204] = 16'h3de0;
mem_array[11207] = 16'h1630;
mem_array[11206] = 16'hbebd;
mem_array[11209] = 16'h8881;
mem_array[11208] = 16'h3e5b;
mem_array[11211] = 16'hecf1;
mem_array[11210] = 16'hbe68;
mem_array[11213] = 16'he9b3;
mem_array[11212] = 16'h3e7d;
mem_array[11215] = 16'hf76b;
mem_array[11214] = 16'hbd8c;
mem_array[11217] = 16'h8fd5;
mem_array[11216] = 16'h3ddd;
mem_array[11219] = 16'ha76c;
mem_array[11218] = 16'hbefb;
mem_array[11221] = 16'h601c;
mem_array[11220] = 16'hbc6e;
mem_array[11223] = 16'h69e2;
mem_array[11222] = 16'h3d1e;
mem_array[11225] = 16'h4b39;
mem_array[11224] = 16'hbe12;
mem_array[11227] = 16'h13fd;
mem_array[11226] = 16'hbe9f;
mem_array[11229] = 16'h4be4;
mem_array[11228] = 16'h3e6d;
mem_array[11231] = 16'h248c;
mem_array[11230] = 16'h3e3e;
mem_array[11233] = 16'hd9d0;
mem_array[11232] = 16'hbe12;
mem_array[11235] = 16'h5821;
mem_array[11234] = 16'h3e32;
mem_array[11237] = 16'h59e2;
mem_array[11236] = 16'h3ef2;
mem_array[11239] = 16'h4aa3;
mem_array[11238] = 16'hbef1;
mem_array[11241] = 16'hcd78;
mem_array[11240] = 16'h3b83;
mem_array[11243] = 16'h1f92;
mem_array[11242] = 16'hbdf7;
mem_array[11245] = 16'h2c8e;
mem_array[11244] = 16'hbe23;
mem_array[11247] = 16'h361f;
mem_array[11246] = 16'hbddc;
mem_array[11249] = 16'hd3d6;
mem_array[11248] = 16'h3e62;
mem_array[11251] = 16'hc6f3;
mem_array[11250] = 16'hbe96;
mem_array[11253] = 16'hf12a;
mem_array[11252] = 16'h3d91;
mem_array[11255] = 16'h70a9;
mem_array[11254] = 16'h3e34;
mem_array[11257] = 16'ha264;
mem_array[11256] = 16'hbe0f;
mem_array[11259] = 16'h99d5;
mem_array[11258] = 16'hbedb;
mem_array[11261] = 16'h1d30;
mem_array[11260] = 16'hbf1e;
mem_array[11263] = 16'hd018;
mem_array[11262] = 16'hbbd7;
mem_array[11265] = 16'h81e4;
mem_array[11264] = 16'h3e6d;
mem_array[11267] = 16'h27be;
mem_array[11266] = 16'hbd82;
mem_array[11269] = 16'h57d6;
mem_array[11268] = 16'hbcda;
mem_array[11271] = 16'h7c0c;
mem_array[11270] = 16'hbd9c;
mem_array[11273] = 16'h0cdb;
mem_array[11272] = 16'h3e56;
mem_array[11275] = 16'hb639;
mem_array[11274] = 16'h3d0f;
mem_array[11277] = 16'h2c48;
mem_array[11276] = 16'h3cff;
mem_array[11279] = 16'h8aa2;
mem_array[11278] = 16'hbd82;
mem_array[11281] = 16'h24ee;
mem_array[11280] = 16'hbe3a;
mem_array[11283] = 16'had30;
mem_array[11282] = 16'hbe1c;
mem_array[11285] = 16'h9c43;
mem_array[11284] = 16'hbf05;
mem_array[11287] = 16'h3b53;
mem_array[11286] = 16'hbeb7;
mem_array[11289] = 16'h35e8;
mem_array[11288] = 16'h3e36;
mem_array[11291] = 16'h030e;
mem_array[11290] = 16'h3d93;
mem_array[11293] = 16'h9052;
mem_array[11292] = 16'hbd9d;
mem_array[11295] = 16'h6e97;
mem_array[11294] = 16'h3e3a;
mem_array[11297] = 16'h9b73;
mem_array[11296] = 16'h3dc2;
mem_array[11299] = 16'hc356;
mem_array[11298] = 16'hbfc6;
mem_array[11301] = 16'hccc5;
mem_array[11300] = 16'hbcfe;
mem_array[11303] = 16'ha160;
mem_array[11302] = 16'hbc80;
mem_array[11305] = 16'he0ce;
mem_array[11304] = 16'hbde3;
mem_array[11307] = 16'hcae8;
mem_array[11306] = 16'hbe99;
mem_array[11309] = 16'h0ab8;
mem_array[11308] = 16'h3e24;
mem_array[11311] = 16'he81d;
mem_array[11310] = 16'hbd95;
mem_array[11313] = 16'h2645;
mem_array[11312] = 16'h3db1;
mem_array[11315] = 16'ha56b;
mem_array[11314] = 16'h3de7;
mem_array[11317] = 16'hf17b;
mem_array[11316] = 16'hbe9b;
mem_array[11319] = 16'h46ba;
mem_array[11318] = 16'h3c1c;
mem_array[11321] = 16'he0e8;
mem_array[11320] = 16'h3dc8;
mem_array[11323] = 16'h73fb;
mem_array[11322] = 16'h3e37;
mem_array[11325] = 16'hd839;
mem_array[11324] = 16'h3ebc;
mem_array[11327] = 16'hd1b2;
mem_array[11326] = 16'hbe33;
mem_array[11329] = 16'h7463;
mem_array[11328] = 16'hbe14;
mem_array[11331] = 16'hebfe;
mem_array[11330] = 16'hbe53;
mem_array[11333] = 16'h0b1b;
mem_array[11332] = 16'h3e87;
mem_array[11335] = 16'h7317;
mem_array[11334] = 16'h3d89;
mem_array[11337] = 16'hecf3;
mem_array[11336] = 16'hbe5a;
mem_array[11339] = 16'h8838;
mem_array[11338] = 16'hbe98;
mem_array[11341] = 16'h5987;
mem_array[11340] = 16'hbe41;
mem_array[11343] = 16'he90c;
mem_array[11342] = 16'h3e15;
mem_array[11345] = 16'hf61f;
mem_array[11344] = 16'h3d57;
mem_array[11347] = 16'hb131;
mem_array[11346] = 16'hbc28;
mem_array[11349] = 16'h5a9a;
mem_array[11348] = 16'hbda6;
mem_array[11351] = 16'h654c;
mem_array[11350] = 16'h3e4a;
mem_array[11353] = 16'h9c8c;
mem_array[11352] = 16'h3e64;
mem_array[11355] = 16'hb2ae;
mem_array[11354] = 16'hbce2;
mem_array[11357] = 16'hb48a;
mem_array[11356] = 16'hbeb3;
mem_array[11359] = 16'h6e1e;
mem_array[11358] = 16'h3dab;
mem_array[11361] = 16'h1fdd;
mem_array[11360] = 16'hbddc;
mem_array[11363] = 16'h585c;
mem_array[11362] = 16'hbc6e;
mem_array[11365] = 16'h3a1d;
mem_array[11364] = 16'h3c1f;
mem_array[11367] = 16'hf0a4;
mem_array[11366] = 16'hbe93;
mem_array[11369] = 16'hed1a;
mem_array[11368] = 16'h3e26;
mem_array[11371] = 16'hf7d0;
mem_array[11370] = 16'hbc82;
mem_array[11373] = 16'h8295;
mem_array[11372] = 16'hbd18;
mem_array[11375] = 16'hc45e;
mem_array[11374] = 16'hbd51;
mem_array[11377] = 16'h0918;
mem_array[11376] = 16'h3e15;
mem_array[11379] = 16'h3d01;
mem_array[11378] = 16'h3cf6;
mem_array[11381] = 16'h23f0;
mem_array[11380] = 16'hbe01;
mem_array[11383] = 16'h09c2;
mem_array[11382] = 16'h3cda;
mem_array[11385] = 16'hd3bb;
mem_array[11384] = 16'hbf34;
mem_array[11387] = 16'hcf36;
mem_array[11386] = 16'hbe51;
mem_array[11389] = 16'habfd;
mem_array[11388] = 16'hbec1;
mem_array[11391] = 16'ha559;
mem_array[11390] = 16'h3daf;
mem_array[11393] = 16'h9e6f;
mem_array[11392] = 16'h3e75;
mem_array[11395] = 16'hc43e;
mem_array[11394] = 16'h3ea4;
mem_array[11397] = 16'h6402;
mem_array[11396] = 16'h3eb4;
mem_array[11399] = 16'hf1f3;
mem_array[11398] = 16'h3e0d;
mem_array[11401] = 16'h1fc5;
mem_array[11400] = 16'h3d5f;
mem_array[11403] = 16'h5e25;
mem_array[11402] = 16'h3eaa;
mem_array[11405] = 16'h4218;
mem_array[11404] = 16'h3ec0;
mem_array[11407] = 16'h7814;
mem_array[11406] = 16'h3ec4;
mem_array[11409] = 16'h4784;
mem_array[11408] = 16'hbe33;
mem_array[11411] = 16'h6567;
mem_array[11410] = 16'h3dc6;
mem_array[11413] = 16'h280d;
mem_array[11412] = 16'hbe9b;
mem_array[11415] = 16'hd5dc;
mem_array[11414] = 16'hbd2d;
mem_array[11417] = 16'he910;
mem_array[11416] = 16'hbf80;
mem_array[11419] = 16'h5e38;
mem_array[11418] = 16'hbf32;
mem_array[11421] = 16'h4b02;
mem_array[11420] = 16'h3d61;
mem_array[11423] = 16'hbaeb;
mem_array[11422] = 16'hbd08;
mem_array[11425] = 16'h6958;
mem_array[11424] = 16'hbe8f;
mem_array[11427] = 16'h701f;
mem_array[11426] = 16'h3e7e;
mem_array[11429] = 16'h82ba;
mem_array[11428] = 16'hbdf2;
mem_array[11431] = 16'h02c8;
mem_array[11430] = 16'hbe51;
mem_array[11433] = 16'h3335;
mem_array[11432] = 16'hbe89;
mem_array[11435] = 16'h6705;
mem_array[11434] = 16'h3e81;
mem_array[11437] = 16'h5b74;
mem_array[11436] = 16'hbec5;
mem_array[11439] = 16'h1869;
mem_array[11438] = 16'h3cfa;
mem_array[11441] = 16'h888c;
mem_array[11440] = 16'h3dc0;
mem_array[11443] = 16'hdeba;
mem_array[11442] = 16'hbd1c;
mem_array[11445] = 16'hba9d;
mem_array[11444] = 16'h3e3f;
mem_array[11447] = 16'hc490;
mem_array[11446] = 16'hbe38;
mem_array[11449] = 16'hd636;
mem_array[11448] = 16'hbe01;
mem_array[11451] = 16'h3251;
mem_array[11450] = 16'hbf4d;
mem_array[11453] = 16'h71ef;
mem_array[11452] = 16'h3d63;
mem_array[11455] = 16'hd48a;
mem_array[11454] = 16'h3ea0;
mem_array[11457] = 16'h25b2;
mem_array[11456] = 16'h3ebb;
mem_array[11459] = 16'hd9ad;
mem_array[11458] = 16'h3e87;
mem_array[11461] = 16'hf7ed;
mem_array[11460] = 16'hbe83;
mem_array[11463] = 16'h0c39;
mem_array[11462] = 16'hbe43;
mem_array[11465] = 16'h8248;
mem_array[11464] = 16'h3c28;
mem_array[11467] = 16'ha9ad;
mem_array[11466] = 16'h3e44;
mem_array[11469] = 16'h8517;
mem_array[11468] = 16'h3da0;
mem_array[11471] = 16'h2a5e;
mem_array[11470] = 16'h3efb;
mem_array[11473] = 16'h81aa;
mem_array[11472] = 16'hbfc7;
mem_array[11475] = 16'hdee1;
mem_array[11474] = 16'hbe14;
mem_array[11477] = 16'h142c;
mem_array[11476] = 16'hbffa;
mem_array[11479] = 16'h6e5e;
mem_array[11478] = 16'hbef2;
mem_array[11481] = 16'h2eb9;
mem_array[11480] = 16'hbd98;
mem_array[11483] = 16'he2bd;
mem_array[11482] = 16'h3daf;
mem_array[11485] = 16'h9159;
mem_array[11484] = 16'hbf71;
mem_array[11487] = 16'hbf28;
mem_array[11486] = 16'hbf07;
mem_array[11489] = 16'hd304;
mem_array[11488] = 16'hbee8;
mem_array[11491] = 16'hfde9;
mem_array[11490] = 16'hbdfd;
mem_array[11493] = 16'hf039;
mem_array[11492] = 16'hbe19;
mem_array[11495] = 16'h43b8;
mem_array[11494] = 16'h3e8b;
mem_array[11497] = 16'hf741;
mem_array[11496] = 16'hbf71;
mem_array[11499] = 16'h8e18;
mem_array[11498] = 16'h3ebb;
mem_array[11501] = 16'ha2b4;
mem_array[11500] = 16'h3ef4;
mem_array[11503] = 16'h8cff;
mem_array[11502] = 16'h3ca4;
mem_array[11505] = 16'h95d1;
mem_array[11504] = 16'hbd02;
mem_array[11507] = 16'hc415;
mem_array[11506] = 16'hbe0e;
mem_array[11509] = 16'h2a68;
mem_array[11508] = 16'hbea9;
mem_array[11511] = 16'h0326;
mem_array[11510] = 16'hbf09;
mem_array[11513] = 16'h8329;
mem_array[11512] = 16'h3e24;
mem_array[11515] = 16'h37ee;
mem_array[11514] = 16'h3da0;
mem_array[11517] = 16'h8969;
mem_array[11516] = 16'hbf5b;
mem_array[11519] = 16'h12db;
mem_array[11518] = 16'h3d7d;
mem_array[11521] = 16'haf76;
mem_array[11520] = 16'hbefd;
mem_array[11523] = 16'h92ac;
mem_array[11522] = 16'h3dca;
mem_array[11525] = 16'ha37d;
mem_array[11524] = 16'hbe5d;
mem_array[11527] = 16'h64a1;
mem_array[11526] = 16'hbf04;
mem_array[11529] = 16'hf1bb;
mem_array[11528] = 16'h3d2a;
mem_array[11531] = 16'hd6c1;
mem_array[11530] = 16'h3eb1;
mem_array[11533] = 16'h7cd8;
mem_array[11532] = 16'hc028;
mem_array[11535] = 16'h60ec;
mem_array[11534] = 16'h3ec7;
mem_array[11537] = 16'h3541;
mem_array[11536] = 16'hbfcd;
mem_array[11539] = 16'hffba;
mem_array[11538] = 16'hbebb;
mem_array[11541] = 16'hfcc1;
mem_array[11540] = 16'hbdbb;
mem_array[11543] = 16'hd6ab;
mem_array[11542] = 16'h3caf;
mem_array[11545] = 16'h3ab6;
mem_array[11544] = 16'hbfac;
mem_array[11547] = 16'ha28a;
mem_array[11546] = 16'hc00d;
mem_array[11549] = 16'h291c;
mem_array[11548] = 16'hbf78;
mem_array[11551] = 16'h74b1;
mem_array[11550] = 16'hbe43;
mem_array[11553] = 16'haab1;
mem_array[11552] = 16'h3e63;
mem_array[11555] = 16'hcf41;
mem_array[11554] = 16'hbf33;
mem_array[11557] = 16'hb867;
mem_array[11556] = 16'hbf04;
mem_array[11559] = 16'h1c6f;
mem_array[11558] = 16'h3ead;
mem_array[11561] = 16'h530f;
mem_array[11560] = 16'h3ea0;
mem_array[11563] = 16'h8084;
mem_array[11562] = 16'hba28;
mem_array[11565] = 16'h4188;
mem_array[11564] = 16'hbd6e;
mem_array[11567] = 16'h6d32;
mem_array[11566] = 16'hbea2;
mem_array[11569] = 16'h8e86;
mem_array[11568] = 16'hbf27;
mem_array[11571] = 16'h4c15;
mem_array[11570] = 16'hbcd2;
mem_array[11573] = 16'h3c1e;
mem_array[11572] = 16'h3ebb;
mem_array[11575] = 16'hebe1;
mem_array[11574] = 16'h3e34;
mem_array[11577] = 16'hd979;
mem_array[11576] = 16'hbf90;
mem_array[11579] = 16'h5922;
mem_array[11578] = 16'hbf1b;
mem_array[11581] = 16'he102;
mem_array[11580] = 16'hbf14;
mem_array[11583] = 16'h1934;
mem_array[11582] = 16'h3e91;
mem_array[11585] = 16'h6f7c;
mem_array[11584] = 16'hbff2;
mem_array[11587] = 16'hd6bd;
mem_array[11586] = 16'hbfe5;
mem_array[11589] = 16'h1769;
mem_array[11588] = 16'hbf9d;
mem_array[11591] = 16'hb720;
mem_array[11590] = 16'h3f61;
mem_array[11593] = 16'hc633;
mem_array[11592] = 16'hbf8c;
mem_array[11595] = 16'h4f45;
mem_array[11594] = 16'hbd89;
mem_array[11597] = 16'haebd;
mem_array[11596] = 16'hbece;
mem_array[11599] = 16'h9f16;
mem_array[11598] = 16'h3eb6;
mem_array[11601] = 16'h2fdd;
mem_array[11600] = 16'h3d3e;
mem_array[11603] = 16'h580d;
mem_array[11602] = 16'h3d84;
mem_array[11605] = 16'h683a;
mem_array[11604] = 16'hbf63;
mem_array[11607] = 16'h9c16;
mem_array[11606] = 16'hbe94;
mem_array[11609] = 16'h2fb8;
mem_array[11608] = 16'hc019;
mem_array[11611] = 16'h493d;
mem_array[11610] = 16'hbe3a;
mem_array[11613] = 16'h4f3d;
mem_array[11612] = 16'hbf39;
mem_array[11615] = 16'h6870;
mem_array[11614] = 16'hbe84;
mem_array[11617] = 16'h8d36;
mem_array[11616] = 16'hbd98;
mem_array[11619] = 16'h8bd6;
mem_array[11618] = 16'h3e87;
mem_array[11621] = 16'h9648;
mem_array[11620] = 16'hbeda;
mem_array[11623] = 16'h9fc1;
mem_array[11622] = 16'h3e31;
mem_array[11625] = 16'h9cf9;
mem_array[11624] = 16'hbf4b;
mem_array[11627] = 16'h1fbd;
mem_array[11626] = 16'h3e8e;
mem_array[11629] = 16'h1925;
mem_array[11628] = 16'hbfa6;
mem_array[11631] = 16'hf6d1;
mem_array[11630] = 16'hbe9b;
mem_array[11633] = 16'h4974;
mem_array[11632] = 16'h3f30;
mem_array[11635] = 16'ha785;
mem_array[11634] = 16'h3e00;
mem_array[11637] = 16'h4292;
mem_array[11636] = 16'hbe98;
mem_array[11639] = 16'h13a8;
mem_array[11638] = 16'hbf1a;
mem_array[11641] = 16'h091e;
mem_array[11640] = 16'hbf01;
mem_array[11643] = 16'h19fe;
mem_array[11642] = 16'hbf1d;
mem_array[11645] = 16'h80a8;
mem_array[11644] = 16'hbdd4;
mem_array[11647] = 16'hfb61;
mem_array[11646] = 16'hbfc5;
mem_array[11649] = 16'hb4e0;
mem_array[11648] = 16'h3e53;
mem_array[11651] = 16'h6cf6;
mem_array[11650] = 16'h3f77;
mem_array[11653] = 16'hca89;
mem_array[11652] = 16'hbe0f;
mem_array[11655] = 16'h31f4;
mem_array[11654] = 16'h3e17;
mem_array[11657] = 16'hb0ca;
mem_array[11656] = 16'h3c2e;
mem_array[11659] = 16'hb3b3;
mem_array[11658] = 16'h3e5c;
mem_array[11661] = 16'h125b;
mem_array[11660] = 16'hbac9;
mem_array[11663] = 16'h075d;
mem_array[11662] = 16'h3d79;
mem_array[11665] = 16'hd0c9;
mem_array[11664] = 16'h3f25;
mem_array[11667] = 16'h153e;
mem_array[11666] = 16'h3e1b;
mem_array[11669] = 16'h0401;
mem_array[11668] = 16'hbe87;
mem_array[11671] = 16'h1fe9;
mem_array[11670] = 16'h3e7d;
mem_array[11673] = 16'hcccc;
mem_array[11672] = 16'hbb0d;
mem_array[11675] = 16'hedb8;
mem_array[11674] = 16'hbdcc;
mem_array[11677] = 16'h48e0;
mem_array[11676] = 16'hbec4;
mem_array[11679] = 16'h2804;
mem_array[11678] = 16'hbc66;
mem_array[11681] = 16'h567f;
mem_array[11680] = 16'h3fd1;
mem_array[11683] = 16'hf8e6;
mem_array[11682] = 16'hbeb6;
mem_array[11685] = 16'h0fe9;
mem_array[11684] = 16'hbf21;
mem_array[11687] = 16'h012c;
mem_array[11686] = 16'hbf5d;
mem_array[11689] = 16'h639e;
mem_array[11688] = 16'hbef2;
mem_array[11691] = 16'h575f;
mem_array[11690] = 16'hbf0c;
mem_array[11693] = 16'hda38;
mem_array[11692] = 16'h3ea1;
mem_array[11695] = 16'h1e9c;
mem_array[11694] = 16'h3ee6;
mem_array[11697] = 16'hd635;
mem_array[11696] = 16'hbd40;
mem_array[11699] = 16'h4476;
mem_array[11698] = 16'hc003;
mem_array[11701] = 16'hc150;
mem_array[11700] = 16'hbf0a;
mem_array[11703] = 16'h39a7;
mem_array[11702] = 16'hbed1;
mem_array[11705] = 16'hb2e2;
mem_array[11704] = 16'h3e90;
mem_array[11707] = 16'h2502;
mem_array[11706] = 16'hbf41;
mem_array[11709] = 16'hf9b0;
mem_array[11708] = 16'hbf6a;
mem_array[11711] = 16'h9fea;
mem_array[11710] = 16'h3ded;
mem_array[11713] = 16'hae13;
mem_array[11712] = 16'h3d4b;
mem_array[11715] = 16'hb5cc;
mem_array[11714] = 16'hbea5;
mem_array[11717] = 16'hfa88;
mem_array[11716] = 16'hbca3;
mem_array[11719] = 16'h9ee5;
mem_array[11718] = 16'h3ec6;
mem_array[11721] = 16'h3892;
mem_array[11720] = 16'h3c86;
mem_array[11723] = 16'hfbc0;
mem_array[11722] = 16'h3b3f;
mem_array[11725] = 16'h679c;
mem_array[11724] = 16'hbe44;
mem_array[11727] = 16'hfe76;
mem_array[11726] = 16'h3e3c;
mem_array[11729] = 16'h259e;
mem_array[11728] = 16'hbe36;
mem_array[11731] = 16'hb747;
mem_array[11730] = 16'h3fa0;
mem_array[11733] = 16'he527;
mem_array[11732] = 16'hbbb6;
mem_array[11735] = 16'h5fa0;
mem_array[11734] = 16'h3e89;
mem_array[11737] = 16'hce83;
mem_array[11736] = 16'hbf59;
mem_array[11739] = 16'h7317;
mem_array[11738] = 16'hbf96;
mem_array[11741] = 16'h82ad;
mem_array[11740] = 16'h3f3e;
mem_array[11743] = 16'h00d4;
mem_array[11742] = 16'h3fba;
mem_array[11745] = 16'h3197;
mem_array[11744] = 16'hbe56;
mem_array[11747] = 16'hdc7f;
mem_array[11746] = 16'h3ed8;
mem_array[11749] = 16'hfda5;
mem_array[11748] = 16'hbec0;
mem_array[11751] = 16'h817a;
mem_array[11750] = 16'h3daa;
mem_array[11753] = 16'h0c8e;
mem_array[11752] = 16'h3e23;
mem_array[11755] = 16'hebfa;
mem_array[11754] = 16'h3f73;
mem_array[11757] = 16'h2821;
mem_array[11756] = 16'h3c35;
mem_array[11759] = 16'h1703;
mem_array[11758] = 16'hbf69;
mem_array[11761] = 16'h9da6;
mem_array[11760] = 16'hbd8d;
mem_array[11763] = 16'h1ae6;
mem_array[11762] = 16'hbc8b;
mem_array[11765] = 16'h925c;
mem_array[11764] = 16'hbc82;
mem_array[11767] = 16'h90cc;
mem_array[11766] = 16'h3cee;
mem_array[11769] = 16'hee7e;
mem_array[11768] = 16'hbc07;
mem_array[11771] = 16'h700b;
mem_array[11770] = 16'hbd0c;
mem_array[11773] = 16'h5f7d;
mem_array[11772] = 16'hbd48;
mem_array[11775] = 16'h6bf9;
mem_array[11774] = 16'h3d9e;
mem_array[11777] = 16'h8f50;
mem_array[11776] = 16'h3dae;
mem_array[11779] = 16'h196e;
mem_array[11778] = 16'hbd09;
mem_array[11781] = 16'h62a3;
mem_array[11780] = 16'hbd1c;
mem_array[11783] = 16'h375a;
mem_array[11782] = 16'hbb94;
mem_array[11785] = 16'hd442;
mem_array[11784] = 16'h3bbc;
mem_array[11787] = 16'hb773;
mem_array[11786] = 16'h3d0e;
mem_array[11789] = 16'h015a;
mem_array[11788] = 16'h3c1e;
mem_array[11791] = 16'h1aa1;
mem_array[11790] = 16'h3c80;
mem_array[11793] = 16'hd517;
mem_array[11792] = 16'h3b5d;
mem_array[11795] = 16'h90e5;
mem_array[11794] = 16'hbd41;
mem_array[11797] = 16'hd107;
mem_array[11796] = 16'h3d7a;
mem_array[11799] = 16'h69ac;
mem_array[11798] = 16'h3d17;
mem_array[11801] = 16'h073d;
mem_array[11800] = 16'hbdac;
mem_array[11803] = 16'h85f6;
mem_array[11802] = 16'hbd9f;
mem_array[11805] = 16'h739d;
mem_array[11804] = 16'hbd22;
mem_array[11807] = 16'h0f37;
mem_array[11806] = 16'hbcbb;
mem_array[11809] = 16'h2441;
mem_array[11808] = 16'h3db0;
mem_array[11811] = 16'h2cd9;
mem_array[11810] = 16'hbdc1;
mem_array[11813] = 16'h50fc;
mem_array[11812] = 16'hbd08;
mem_array[11815] = 16'hdca5;
mem_array[11814] = 16'hbcfe;
mem_array[11817] = 16'h9436;
mem_array[11816] = 16'h3d03;
mem_array[11819] = 16'hd041;
mem_array[11818] = 16'h3d64;
mem_array[11821] = 16'hfa79;
mem_array[11820] = 16'hbca9;
mem_array[11823] = 16'h4c19;
mem_array[11822] = 16'h3ee6;
mem_array[11825] = 16'h5b02;
mem_array[11824] = 16'h3e7e;
mem_array[11827] = 16'hef0c;
mem_array[11826] = 16'h3db9;
mem_array[11829] = 16'hc185;
mem_array[11828] = 16'h3ea6;
mem_array[11831] = 16'h37be;
mem_array[11830] = 16'hbd88;
mem_array[11833] = 16'h79eb;
mem_array[11832] = 16'h3fbf;
mem_array[11835] = 16'hb4e8;
mem_array[11834] = 16'h3fd7;
mem_array[11837] = 16'hcc33;
mem_array[11836] = 16'h3d50;
mem_array[11839] = 16'hdbfb;
mem_array[11838] = 16'hbd41;
mem_array[11841] = 16'h502a;
mem_array[11840] = 16'h3cca;
mem_array[11843] = 16'h4bc6;
mem_array[11842] = 16'hbd6e;
mem_array[11845] = 16'hd8d7;
mem_array[11844] = 16'hbf17;
mem_array[11847] = 16'hc4c1;
mem_array[11846] = 16'h3de4;
mem_array[11849] = 16'h6643;
mem_array[11848] = 16'hbd4c;
mem_array[11851] = 16'h5216;
mem_array[11850] = 16'hbfa6;
mem_array[11853] = 16'hf9df;
mem_array[11852] = 16'hbd43;
mem_array[11855] = 16'hc777;
mem_array[11854] = 16'hbdc3;
mem_array[11857] = 16'h92e2;
mem_array[11856] = 16'h3dd0;
mem_array[11859] = 16'hb8cf;
mem_array[11858] = 16'h3e5c;
mem_array[11861] = 16'h0214;
mem_array[11860] = 16'hbeee;
mem_array[11863] = 16'he808;
mem_array[11862] = 16'h3e21;
mem_array[11865] = 16'hfb00;
mem_array[11864] = 16'hbd9f;
mem_array[11867] = 16'h5a3e;
mem_array[11866] = 16'hbfe8;
mem_array[11869] = 16'hdb79;
mem_array[11868] = 16'h3fab;
mem_array[11871] = 16'h7f7f;
mem_array[11870] = 16'h3fd4;
mem_array[11873] = 16'h77ef;
mem_array[11872] = 16'h3f0a;
mem_array[11875] = 16'hb274;
mem_array[11874] = 16'h3e84;
mem_array[11877] = 16'h6d01;
mem_array[11876] = 16'h3d12;
mem_array[11879] = 16'h82a6;
mem_array[11878] = 16'hbef6;
mem_array[11881] = 16'h8333;
mem_array[11880] = 16'h3d88;
mem_array[11883] = 16'hc2ec;
mem_array[11882] = 16'h3f1a;
mem_array[11885] = 16'h3015;
mem_array[11884] = 16'hbdb0;
mem_array[11887] = 16'hf8de;
mem_array[11886] = 16'hbf09;
mem_array[11889] = 16'hadf1;
mem_array[11888] = 16'h3eb4;
mem_array[11891] = 16'h7cec;
mem_array[11890] = 16'h3ed1;
mem_array[11893] = 16'h5eba;
mem_array[11892] = 16'hbe67;
mem_array[11895] = 16'h15cd;
mem_array[11894] = 16'h3e87;
mem_array[11897] = 16'he31d;
mem_array[11896] = 16'hbdd0;
mem_array[11899] = 16'h031f;
mem_array[11898] = 16'h3f2d;
mem_array[11901] = 16'hdac6;
mem_array[11900] = 16'h3c38;
mem_array[11903] = 16'h278b;
mem_array[11902] = 16'h3de6;
mem_array[11905] = 16'h14e9;
mem_array[11904] = 16'h3fbe;
mem_array[11907] = 16'h0847;
mem_array[11906] = 16'h4008;
mem_array[11909] = 16'hb7b9;
mem_array[11908] = 16'h3fba;
mem_array[11911] = 16'h5307;
mem_array[11910] = 16'hbf15;
mem_array[11913] = 16'h6cfc;
mem_array[11912] = 16'h3e0d;
mem_array[11915] = 16'h17fa;
mem_array[11914] = 16'hbe3a;
mem_array[11917] = 16'h5f69;
mem_array[11916] = 16'h3ed4;
mem_array[11919] = 16'h723b;
mem_array[11918] = 16'h3f3c;
mem_array[11921] = 16'he974;
mem_array[11920] = 16'h3db1;
mem_array[11923] = 16'h0d43;
mem_array[11922] = 16'hbd9e;
mem_array[11925] = 16'he843;
mem_array[11924] = 16'h3d5b;
mem_array[11927] = 16'h2d30;
mem_array[11926] = 16'hbf6b;
mem_array[11929] = 16'h2977;
mem_array[11928] = 16'hbe8e;
mem_array[11931] = 16'h8cf0;
mem_array[11930] = 16'h3f62;
mem_array[11933] = 16'h92f6;
mem_array[11932] = 16'hbe70;
mem_array[11935] = 16'h5c74;
mem_array[11934] = 16'h3ed7;
mem_array[11937] = 16'hf8f5;
mem_array[11936] = 16'h3f27;
mem_array[11939] = 16'h528e;
mem_array[11938] = 16'hbed7;
mem_array[11941] = 16'h159f;
mem_array[11940] = 16'h3f0d;
mem_array[11943] = 16'h6866;
mem_array[11942] = 16'h3f73;
mem_array[11945] = 16'hd0fa;
mem_array[11944] = 16'h3f4e;
mem_array[11947] = 16'ha91e;
mem_array[11946] = 16'hbf17;
mem_array[11949] = 16'h393d;
mem_array[11948] = 16'h3f30;
mem_array[11951] = 16'h9346;
mem_array[11950] = 16'hbb10;
mem_array[11953] = 16'h0ec3;
mem_array[11952] = 16'h3f37;
mem_array[11955] = 16'h13e7;
mem_array[11954] = 16'h3f86;
mem_array[11957] = 16'ha450;
mem_array[11956] = 16'h3f22;
mem_array[11959] = 16'h8985;
mem_array[11958] = 16'h3ebf;
mem_array[11961] = 16'h80ec;
mem_array[11960] = 16'h3ccf;
mem_array[11963] = 16'h7825;
mem_array[11962] = 16'hbac6;
mem_array[11965] = 16'h22ac;
mem_array[11964] = 16'h3da9;
mem_array[11967] = 16'hdc17;
mem_array[11966] = 16'hbf7a;
mem_array[11969] = 16'hc80a;
mem_array[11968] = 16'hbebc;
mem_array[11971] = 16'hdeae;
mem_array[11970] = 16'hbe79;
mem_array[11973] = 16'h5626;
mem_array[11972] = 16'hbf46;
mem_array[11975] = 16'h4f3d;
mem_array[11974] = 16'h3dc0;
mem_array[11977] = 16'h44c4;
mem_array[11976] = 16'h3fa7;
mem_array[11979] = 16'h2540;
mem_array[11978] = 16'h3cfa;
mem_array[11981] = 16'h4d3d;
mem_array[11980] = 16'h3e05;
mem_array[11983] = 16'hb72d;
mem_array[11982] = 16'h3e38;
mem_array[11985] = 16'h27e7;
mem_array[11984] = 16'hbb84;
mem_array[11987] = 16'h3d59;
mem_array[11986] = 16'hbf88;
mem_array[11989] = 16'hd944;
mem_array[11988] = 16'hbf0e;
mem_array[11991] = 16'h70ff;
mem_array[11990] = 16'h4007;
mem_array[11993] = 16'hf8b1;
mem_array[11992] = 16'h3eeb;
mem_array[11995] = 16'h8114;
mem_array[11994] = 16'h3f19;
mem_array[11997] = 16'h6ec8;
mem_array[11996] = 16'h3eb7;
mem_array[11999] = 16'h5e31;
mem_array[11998] = 16'hbe58;
mem_array[12001] = 16'h72b5;
mem_array[12000] = 16'h3f24;
mem_array[12003] = 16'he354;
mem_array[12002] = 16'h3d8d;
mem_array[12005] = 16'h9a74;
mem_array[12004] = 16'h3df7;
mem_array[12007] = 16'hd958;
mem_array[12006] = 16'h3eec;
mem_array[12009] = 16'h17bb;
mem_array[12008] = 16'hbe8b;
mem_array[12011] = 16'he915;
mem_array[12010] = 16'hbf67;
mem_array[12013] = 16'hb25e;
mem_array[12012] = 16'h3f0d;
mem_array[12015] = 16'hd43d;
mem_array[12014] = 16'h3f0a;
mem_array[12017] = 16'he123;
mem_array[12016] = 16'h3f09;
mem_array[12019] = 16'hac64;
mem_array[12018] = 16'hbe17;
mem_array[12021] = 16'h33f8;
mem_array[12020] = 16'hbb40;
mem_array[12023] = 16'h605d;
mem_array[12022] = 16'h3d4f;
mem_array[12025] = 16'h30f4;
mem_array[12024] = 16'hbf80;
mem_array[12027] = 16'h41c6;
mem_array[12026] = 16'h3ed0;
mem_array[12029] = 16'h89cf;
mem_array[12028] = 16'h3ec4;
mem_array[12031] = 16'h086c;
mem_array[12030] = 16'h3e64;
mem_array[12033] = 16'h9e3b;
mem_array[12032] = 16'hbeab;
mem_array[12035] = 16'h5dcb;
mem_array[12034] = 16'hbed1;
mem_array[12037] = 16'h5668;
mem_array[12036] = 16'hbee3;
mem_array[12039] = 16'h6842;
mem_array[12038] = 16'hbd68;
mem_array[12041] = 16'h61a4;
mem_array[12040] = 16'h3f09;
mem_array[12043] = 16'h7a82;
mem_array[12042] = 16'h3e7a;
mem_array[12045] = 16'h3516;
mem_array[12044] = 16'hbe8e;
mem_array[12047] = 16'h3b29;
mem_array[12046] = 16'hbec7;
mem_array[12049] = 16'h1adf;
mem_array[12048] = 16'hbf04;
mem_array[12051] = 16'h3459;
mem_array[12050] = 16'h3e3d;
mem_array[12053] = 16'hbe73;
mem_array[12052] = 16'h3f1e;
mem_array[12055] = 16'hbbc8;
mem_array[12054] = 16'h3d0e;
mem_array[12057] = 16'h624c;
mem_array[12056] = 16'hbd36;
mem_array[12059] = 16'heb85;
mem_array[12058] = 16'h3f4a;
mem_array[12061] = 16'h6c6f;
mem_array[12060] = 16'h3e09;
mem_array[12063] = 16'hc0a6;
mem_array[12062] = 16'hbe83;
mem_array[12065] = 16'h5f55;
mem_array[12064] = 16'hba45;
mem_array[12067] = 16'he526;
mem_array[12066] = 16'h3efc;
mem_array[12069] = 16'h1fbc;
mem_array[12068] = 16'hbeec;
mem_array[12071] = 16'h2644;
mem_array[12070] = 16'hbf0a;
mem_array[12073] = 16'h5439;
mem_array[12072] = 16'h3eb3;
mem_array[12075] = 16'hdc9f;
mem_array[12074] = 16'h3d92;
mem_array[12077] = 16'h90bb;
mem_array[12076] = 16'h3d86;
mem_array[12079] = 16'hdb1c;
mem_array[12078] = 16'hbf7d;
mem_array[12081] = 16'h4b28;
mem_array[12080] = 16'hbd90;
mem_array[12083] = 16'h7a58;
mem_array[12082] = 16'hbd72;
mem_array[12085] = 16'ha722;
mem_array[12084] = 16'hbf1f;
mem_array[12087] = 16'hba53;
mem_array[12086] = 16'hbe15;
mem_array[12089] = 16'hf89e;
mem_array[12088] = 16'h3f15;
mem_array[12091] = 16'hc689;
mem_array[12090] = 16'hbe39;
mem_array[12093] = 16'h2eca;
mem_array[12092] = 16'hbea9;
mem_array[12095] = 16'h6dc5;
mem_array[12094] = 16'h3e89;
mem_array[12097] = 16'h81de;
mem_array[12096] = 16'hbe25;
mem_array[12099] = 16'hd715;
mem_array[12098] = 16'h3e99;
mem_array[12101] = 16'h3503;
mem_array[12100] = 16'h3ed6;
mem_array[12103] = 16'hd2ce;
mem_array[12102] = 16'h3eab;
mem_array[12105] = 16'hca3e;
mem_array[12104] = 16'hbf00;
mem_array[12107] = 16'hbff7;
mem_array[12106] = 16'hbd74;
mem_array[12109] = 16'ha1cf;
mem_array[12108] = 16'hbe1d;
mem_array[12111] = 16'he05f;
mem_array[12110] = 16'h3d30;
mem_array[12113] = 16'hbb64;
mem_array[12112] = 16'hbe4b;
mem_array[12115] = 16'h3fe3;
mem_array[12114] = 16'hbf24;
mem_array[12117] = 16'hf4c6;
mem_array[12116] = 16'h3eb3;
mem_array[12119] = 16'h82a3;
mem_array[12118] = 16'h3e95;
mem_array[12121] = 16'h61ca;
mem_array[12120] = 16'h3d32;
mem_array[12123] = 16'h1c97;
mem_array[12122] = 16'h3e93;
mem_array[12125] = 16'h1ea2;
mem_array[12124] = 16'h3de8;
mem_array[12127] = 16'ha03e;
mem_array[12126] = 16'h3e98;
mem_array[12129] = 16'h52cb;
mem_array[12128] = 16'hbdb1;
mem_array[12131] = 16'hea5b;
mem_array[12130] = 16'hbc84;
mem_array[12133] = 16'hcd37;
mem_array[12132] = 16'hbd8d;
mem_array[12135] = 16'hd6a7;
mem_array[12134] = 16'hbecb;
mem_array[12137] = 16'h75d9;
mem_array[12136] = 16'h3e64;
mem_array[12139] = 16'h3c8f;
mem_array[12138] = 16'hbec3;
mem_array[12141] = 16'h5ba4;
mem_array[12140] = 16'hbd31;
mem_array[12143] = 16'h83f5;
mem_array[12142] = 16'hbc92;
mem_array[12145] = 16'ha3cd;
mem_array[12144] = 16'hbe36;
mem_array[12147] = 16'hf336;
mem_array[12146] = 16'h3e94;
mem_array[12149] = 16'hccd9;
mem_array[12148] = 16'hbebe;
mem_array[12151] = 16'h4cfd;
mem_array[12150] = 16'hbd5a;
mem_array[12153] = 16'he05b;
mem_array[12152] = 16'hbe8c;
mem_array[12155] = 16'h0627;
mem_array[12154] = 16'h3eb1;
mem_array[12157] = 16'hde38;
mem_array[12156] = 16'h3f15;
mem_array[12159] = 16'h39cf;
mem_array[12158] = 16'h3d85;
mem_array[12161] = 16'h2e58;
mem_array[12160] = 16'hbe85;
mem_array[12163] = 16'h73b5;
mem_array[12162] = 16'h3ac8;
mem_array[12165] = 16'h9d13;
mem_array[12164] = 16'hbf8c;
mem_array[12167] = 16'h0d1c;
mem_array[12166] = 16'hbead;
mem_array[12169] = 16'hed17;
mem_array[12168] = 16'h3d1d;
mem_array[12171] = 16'h11d9;
mem_array[12170] = 16'h3f08;
mem_array[12173] = 16'h948b;
mem_array[12172] = 16'hbe99;
mem_array[12175] = 16'h3352;
mem_array[12174] = 16'hbe07;
mem_array[12177] = 16'h6807;
mem_array[12176] = 16'h3f45;
mem_array[12179] = 16'h0dfd;
mem_array[12178] = 16'hbd03;
mem_array[12181] = 16'h363b;
mem_array[12180] = 16'h3e12;
mem_array[12183] = 16'hf5d8;
mem_array[12182] = 16'h3f68;
mem_array[12185] = 16'h4b06;
mem_array[12184] = 16'h3db3;
mem_array[12187] = 16'h6a6b;
mem_array[12186] = 16'h3e17;
mem_array[12189] = 16'h41f4;
mem_array[12188] = 16'h3ccc;
mem_array[12191] = 16'h49ed;
mem_array[12190] = 16'hbeff;
mem_array[12193] = 16'h1868;
mem_array[12192] = 16'h3e15;
mem_array[12195] = 16'h73d8;
mem_array[12194] = 16'hbea9;
mem_array[12197] = 16'h0756;
mem_array[12196] = 16'h3e65;
mem_array[12199] = 16'h2256;
mem_array[12198] = 16'h3e59;
mem_array[12201] = 16'h5eba;
mem_array[12200] = 16'h3d89;
mem_array[12203] = 16'ha199;
mem_array[12202] = 16'h3d2c;
mem_array[12205] = 16'hfbf7;
mem_array[12204] = 16'hbb46;
mem_array[12207] = 16'h8ce4;
mem_array[12206] = 16'h3e7d;
mem_array[12209] = 16'hd8c1;
mem_array[12208] = 16'hbe60;
mem_array[12211] = 16'h3cc0;
mem_array[12210] = 16'hbdc8;
mem_array[12213] = 16'h44c4;
mem_array[12212] = 16'h3d1f;
mem_array[12215] = 16'h5496;
mem_array[12214] = 16'h3d37;
mem_array[12217] = 16'haeaa;
mem_array[12216] = 16'h3bdf;
mem_array[12219] = 16'h47cd;
mem_array[12218] = 16'h3d50;
mem_array[12221] = 16'hde0a;
mem_array[12220] = 16'hbf03;
mem_array[12223] = 16'hbe63;
mem_array[12222] = 16'hbc89;
mem_array[12225] = 16'h348c;
mem_array[12224] = 16'hbe55;
mem_array[12227] = 16'h08d7;
mem_array[12226] = 16'hbc81;
mem_array[12229] = 16'ha6ea;
mem_array[12228] = 16'hbd6f;
mem_array[12231] = 16'h94fa;
mem_array[12230] = 16'h3ec0;
mem_array[12233] = 16'hfb37;
mem_array[12232] = 16'hbe3c;
mem_array[12235] = 16'h7619;
mem_array[12234] = 16'h3f1c;
mem_array[12237] = 16'h768f;
mem_array[12236] = 16'h3f0a;
mem_array[12239] = 16'hd3ea;
mem_array[12238] = 16'hbd80;
mem_array[12241] = 16'h740a;
mem_array[12240] = 16'h3dd6;
mem_array[12243] = 16'ha425;
mem_array[12242] = 16'h3e64;
mem_array[12245] = 16'h4346;
mem_array[12244] = 16'hbe5f;
mem_array[12247] = 16'haa6b;
mem_array[12246] = 16'hbf02;
mem_array[12249] = 16'h2415;
mem_array[12248] = 16'hbe90;
mem_array[12251] = 16'h1fb4;
mem_array[12250] = 16'hbeaa;
mem_array[12253] = 16'hf635;
mem_array[12252] = 16'h3c81;
mem_array[12255] = 16'hb86f;
mem_array[12254] = 16'hbedd;
mem_array[12257] = 16'hddfc;
mem_array[12256] = 16'h3e04;
mem_array[12259] = 16'h27c7;
mem_array[12258] = 16'hbe15;
mem_array[12261] = 16'h2cc8;
mem_array[12260] = 16'hbd24;
mem_array[12263] = 16'h6dae;
mem_array[12262] = 16'h3c41;
mem_array[12265] = 16'heb5c;
mem_array[12264] = 16'hbe27;
mem_array[12267] = 16'h4ca0;
mem_array[12266] = 16'h3e3d;
mem_array[12269] = 16'h026a;
mem_array[12268] = 16'h3d09;
mem_array[12271] = 16'h02d9;
mem_array[12270] = 16'hbe08;
mem_array[12273] = 16'h62a6;
mem_array[12272] = 16'h3e6d;
mem_array[12275] = 16'h13ea;
mem_array[12274] = 16'h3de7;
mem_array[12277] = 16'hf09b;
mem_array[12276] = 16'hbecc;
mem_array[12279] = 16'h7698;
mem_array[12278] = 16'h3e27;
mem_array[12281] = 16'h5959;
mem_array[12280] = 16'h3e3a;
mem_array[12283] = 16'ha876;
mem_array[12282] = 16'h3d98;
mem_array[12285] = 16'h656f;
mem_array[12284] = 16'hbeff;
mem_array[12287] = 16'heb38;
mem_array[12286] = 16'hbe25;
mem_array[12289] = 16'h0d4f;
mem_array[12288] = 16'h3dfd;
mem_array[12291] = 16'h7307;
mem_array[12290] = 16'hbdbc;
mem_array[12293] = 16'hb88e;
mem_array[12292] = 16'h3ec9;
mem_array[12295] = 16'h892d;
mem_array[12294] = 16'h3d77;
mem_array[12297] = 16'h1d3b;
mem_array[12296] = 16'h3eaa;
mem_array[12299] = 16'he1ec;
mem_array[12298] = 16'hbe91;
mem_array[12301] = 16'hc941;
mem_array[12300] = 16'h3ecd;
mem_array[12303] = 16'h32f6;
mem_array[12302] = 16'hbd37;
mem_array[12305] = 16'h1dfc;
mem_array[12304] = 16'h3d8b;
mem_array[12307] = 16'h4224;
mem_array[12306] = 16'hbe01;
mem_array[12309] = 16'h00ee;
mem_array[12308] = 16'hbea3;
mem_array[12311] = 16'hfe47;
mem_array[12310] = 16'h3ddb;
mem_array[12313] = 16'hcce6;
mem_array[12312] = 16'h3d7b;
mem_array[12315] = 16'h48c9;
mem_array[12314] = 16'hbeb0;
mem_array[12317] = 16'h1f3f;
mem_array[12316] = 16'hbc4a;
mem_array[12319] = 16'h3b64;
mem_array[12318] = 16'h3e4d;
mem_array[12321] = 16'h3f36;
mem_array[12320] = 16'hbb13;
mem_array[12323] = 16'h8591;
mem_array[12322] = 16'hbd41;
mem_array[12325] = 16'h1b5a;
mem_array[12324] = 16'hbe88;
mem_array[12327] = 16'h6f16;
mem_array[12326] = 16'h3e29;
mem_array[12329] = 16'hd495;
mem_array[12328] = 16'h3e21;
mem_array[12331] = 16'h22b8;
mem_array[12330] = 16'hbe5f;
mem_array[12333] = 16'hb74b;
mem_array[12332] = 16'hbd5a;
mem_array[12335] = 16'hd634;
mem_array[12334] = 16'hbe80;
mem_array[12337] = 16'h90d4;
mem_array[12336] = 16'hbded;
mem_array[12339] = 16'h5904;
mem_array[12338] = 16'h3cc2;
mem_array[12341] = 16'hb216;
mem_array[12340] = 16'h3ebf;
mem_array[12343] = 16'hfb9c;
mem_array[12342] = 16'hbe02;
mem_array[12345] = 16'h26f6;
mem_array[12344] = 16'hbd8f;
mem_array[12347] = 16'ha177;
mem_array[12346] = 16'hbe80;
mem_array[12349] = 16'h681a;
mem_array[12348] = 16'h3ee8;
mem_array[12351] = 16'h1853;
mem_array[12350] = 16'h3f43;
mem_array[12353] = 16'had7d;
mem_array[12352] = 16'h3e08;
mem_array[12355] = 16'h5852;
mem_array[12354] = 16'hbe59;
mem_array[12357] = 16'heade;
mem_array[12356] = 16'h3e09;
mem_array[12359] = 16'hd949;
mem_array[12358] = 16'hbf5a;
mem_array[12361] = 16'hbe98;
mem_array[12360] = 16'hbe76;
mem_array[12363] = 16'ha994;
mem_array[12362] = 16'hbeae;
mem_array[12365] = 16'hcb6b;
mem_array[12364] = 16'h3d04;
mem_array[12367] = 16'h4381;
mem_array[12366] = 16'h3ea2;
mem_array[12369] = 16'hd8bc;
mem_array[12368] = 16'h3d20;
mem_array[12371] = 16'hbef5;
mem_array[12370] = 16'h3efe;
mem_array[12373] = 16'hc841;
mem_array[12372] = 16'hbddc;
mem_array[12375] = 16'h0a1c;
mem_array[12374] = 16'hbd9f;
mem_array[12377] = 16'h5b82;
mem_array[12376] = 16'hbe91;
mem_array[12379] = 16'h4bf0;
mem_array[12378] = 16'hbe36;
mem_array[12381] = 16'h9a2c;
mem_array[12380] = 16'hbd86;
mem_array[12383] = 16'h2e41;
mem_array[12382] = 16'hbd8e;
mem_array[12385] = 16'h973c;
mem_array[12384] = 16'h3c18;
mem_array[12387] = 16'hf45b;
mem_array[12386] = 16'h3ddd;
mem_array[12389] = 16'h5891;
mem_array[12388] = 16'h3cc8;
mem_array[12391] = 16'h4d26;
mem_array[12390] = 16'hbc12;
mem_array[12393] = 16'h9ed8;
mem_array[12392] = 16'h3b16;
mem_array[12395] = 16'hfb30;
mem_array[12394] = 16'h3ada;
mem_array[12397] = 16'hef78;
mem_array[12396] = 16'h3dd9;
mem_array[12399] = 16'h4e57;
mem_array[12398] = 16'hbe72;
mem_array[12401] = 16'h118e;
mem_array[12400] = 16'hbe88;
mem_array[12403] = 16'h73d4;
mem_array[12402] = 16'hbde0;
mem_array[12405] = 16'h3b89;
mem_array[12404] = 16'hbf42;
mem_array[12407] = 16'hcb96;
mem_array[12406] = 16'hbe22;
mem_array[12409] = 16'h1edf;
mem_array[12408] = 16'hbd6e;
mem_array[12411] = 16'h406b;
mem_array[12410] = 16'h3f06;
mem_array[12413] = 16'h927d;
mem_array[12412] = 16'hbe65;
mem_array[12415] = 16'h2624;
mem_array[12414] = 16'hbd97;
mem_array[12417] = 16'hb9d7;
mem_array[12416] = 16'h3cbe;
mem_array[12419] = 16'had71;
mem_array[12418] = 16'hbf34;
mem_array[12421] = 16'h3fa9;
mem_array[12420] = 16'hbe77;
mem_array[12423] = 16'h0aed;
mem_array[12422] = 16'hbec5;
mem_array[12425] = 16'hf9df;
mem_array[12424] = 16'hbdf6;
mem_array[12427] = 16'h97d1;
mem_array[12426] = 16'h3e82;
mem_array[12429] = 16'h7ced;
mem_array[12428] = 16'h3ea9;
mem_array[12431] = 16'hccae;
mem_array[12430] = 16'h3e5c;
mem_array[12433] = 16'h3bf1;
mem_array[12432] = 16'hbd9d;
mem_array[12435] = 16'h5a4a;
mem_array[12434] = 16'hbf07;
mem_array[12437] = 16'h8f8b;
mem_array[12436] = 16'hbd4d;
mem_array[12439] = 16'h52a4;
mem_array[12438] = 16'h3c84;
mem_array[12441] = 16'h9bac;
mem_array[12440] = 16'hbba6;
mem_array[12443] = 16'hfd1a;
mem_array[12442] = 16'hbdad;
mem_array[12445] = 16'h4f19;
mem_array[12444] = 16'h3e62;
mem_array[12447] = 16'h60f3;
mem_array[12446] = 16'h3ec1;
mem_array[12449] = 16'h2736;
mem_array[12448] = 16'h3dab;
mem_array[12451] = 16'h5ae3;
mem_array[12450] = 16'h3d77;
mem_array[12453] = 16'he39a;
mem_array[12452] = 16'h3c70;
mem_array[12455] = 16'h7974;
mem_array[12454] = 16'h3e14;
mem_array[12457] = 16'h9584;
mem_array[12456] = 16'h3d8a;
mem_array[12459] = 16'h38e3;
mem_array[12458] = 16'hbe2e;
mem_array[12461] = 16'h68f8;
mem_array[12460] = 16'hbe90;
mem_array[12463] = 16'h668b;
mem_array[12462] = 16'hbdeb;
mem_array[12465] = 16'hc097;
mem_array[12464] = 16'hbeec;
mem_array[12467] = 16'ha0fe;
mem_array[12466] = 16'h3df4;
mem_array[12469] = 16'h5dc2;
mem_array[12468] = 16'h3eb2;
mem_array[12471] = 16'h6d7a;
mem_array[12470] = 16'h3e22;
mem_array[12473] = 16'h7ef6;
mem_array[12472] = 16'hbe02;
mem_array[12475] = 16'h77d0;
mem_array[12474] = 16'hbe38;
mem_array[12477] = 16'h0f31;
mem_array[12476] = 16'h3d71;
mem_array[12479] = 16'hc77a;
mem_array[12478] = 16'hbf07;
mem_array[12481] = 16'h2844;
mem_array[12480] = 16'hbeaf;
mem_array[12483] = 16'h87b9;
mem_array[12482] = 16'hbf11;
mem_array[12485] = 16'h215d;
mem_array[12484] = 16'hbded;
mem_array[12487] = 16'he6cf;
mem_array[12486] = 16'hbd92;
mem_array[12489] = 16'h57cf;
mem_array[12488] = 16'h3e36;
mem_array[12491] = 16'ha4cd;
mem_array[12490] = 16'h3ddb;
mem_array[12493] = 16'h511d;
mem_array[12492] = 16'h3e15;
mem_array[12495] = 16'hfc06;
mem_array[12494] = 16'hbe5d;
mem_array[12497] = 16'hb2ac;
mem_array[12496] = 16'hbda0;
mem_array[12499] = 16'h505e;
mem_array[12498] = 16'h3eda;
mem_array[12501] = 16'hd3f1;
mem_array[12500] = 16'h3d94;
mem_array[12503] = 16'h8f4a;
mem_array[12502] = 16'hbadf;
mem_array[12505] = 16'h35f7;
mem_array[12504] = 16'hbe77;
mem_array[12507] = 16'h4364;
mem_array[12506] = 16'hbdaf;
mem_array[12509] = 16'h7d53;
mem_array[12508] = 16'h3d86;
mem_array[12511] = 16'h1293;
mem_array[12510] = 16'h3dbb;
mem_array[12513] = 16'h786d;
mem_array[12512] = 16'h3e37;
mem_array[12515] = 16'h29c6;
mem_array[12514] = 16'hbd77;
mem_array[12517] = 16'hc8a1;
mem_array[12516] = 16'h3e50;
mem_array[12519] = 16'h7f9e;
mem_array[12518] = 16'hbecc;
mem_array[12521] = 16'hc9c3;
mem_array[12520] = 16'hbf04;
mem_array[12523] = 16'h5f64;
mem_array[12522] = 16'h3bd1;
mem_array[12525] = 16'h93d3;
mem_array[12524] = 16'hbf12;
mem_array[12527] = 16'h9a16;
mem_array[12526] = 16'hbda4;
mem_array[12529] = 16'hbf92;
mem_array[12528] = 16'h3e15;
mem_array[12531] = 16'h2c45;
mem_array[12530] = 16'hbe1e;
mem_array[12533] = 16'h3f2a;
mem_array[12532] = 16'h3d36;
mem_array[12535] = 16'hb2b1;
mem_array[12534] = 16'h3e56;
mem_array[12537] = 16'hf07c;
mem_array[12536] = 16'hbe70;
mem_array[12539] = 16'h1cee;
mem_array[12538] = 16'hbece;
mem_array[12541] = 16'h0ff8;
mem_array[12540] = 16'hbe8e;
mem_array[12543] = 16'hcb0e;
mem_array[12542] = 16'hbedc;
mem_array[12545] = 16'h224f;
mem_array[12544] = 16'hbd5a;
mem_array[12547] = 16'hc56c;
mem_array[12546] = 16'h3c4b;
mem_array[12549] = 16'h279f;
mem_array[12548] = 16'h3e34;
mem_array[12551] = 16'h4047;
mem_array[12550] = 16'hbe90;
mem_array[12553] = 16'h43a3;
mem_array[12552] = 16'h3e8a;
mem_array[12555] = 16'he44f;
mem_array[12554] = 16'hbe37;
mem_array[12557] = 16'hc4d9;
mem_array[12556] = 16'h3e3a;
mem_array[12559] = 16'hfa4d;
mem_array[12558] = 16'hbe72;
mem_array[12561] = 16'hf35f;
mem_array[12560] = 16'hbd9f;
mem_array[12563] = 16'h1708;
mem_array[12562] = 16'hbda2;
mem_array[12565] = 16'hb068;
mem_array[12564] = 16'hbe26;
mem_array[12567] = 16'he337;
mem_array[12566] = 16'h3e91;
mem_array[12569] = 16'h9780;
mem_array[12568] = 16'h3c39;
mem_array[12571] = 16'hf3db;
mem_array[12570] = 16'hbb15;
mem_array[12573] = 16'h7813;
mem_array[12572] = 16'h3e10;
mem_array[12575] = 16'h3d30;
mem_array[12574] = 16'hbd25;
mem_array[12577] = 16'hfa63;
mem_array[12576] = 16'h3e18;
mem_array[12579] = 16'h2924;
mem_array[12578] = 16'h3c98;
mem_array[12581] = 16'h6ba7;
mem_array[12580] = 16'h3c8e;
mem_array[12583] = 16'h9535;
mem_array[12582] = 16'h3e58;
mem_array[12585] = 16'h9a58;
mem_array[12584] = 16'hbee5;
mem_array[12587] = 16'hbd82;
mem_array[12586] = 16'hbe05;
mem_array[12589] = 16'hca1d;
mem_array[12588] = 16'h3e8e;
mem_array[12591] = 16'h5338;
mem_array[12590] = 16'hbe76;
mem_array[12593] = 16'h525a;
mem_array[12592] = 16'hbd8a;
mem_array[12595] = 16'h193a;
mem_array[12594] = 16'hbcad;
mem_array[12597] = 16'hd66d;
mem_array[12596] = 16'hbe2d;
mem_array[12599] = 16'h3fc7;
mem_array[12598] = 16'hbbd0;
mem_array[12601] = 16'hb739;
mem_array[12600] = 16'h3c96;
mem_array[12603] = 16'h96ca;
mem_array[12602] = 16'hbe6e;
mem_array[12605] = 16'h9071;
mem_array[12604] = 16'h3d9e;
mem_array[12607] = 16'hf5b0;
mem_array[12606] = 16'hbd8d;
mem_array[12609] = 16'h62c1;
mem_array[12608] = 16'hbe53;
mem_array[12611] = 16'hea5f;
mem_array[12610] = 16'hbd6c;
mem_array[12613] = 16'h6008;
mem_array[12612] = 16'h3e2f;
mem_array[12615] = 16'h3cf1;
mem_array[12614] = 16'hbda2;
mem_array[12617] = 16'he16b;
mem_array[12616] = 16'hbd3b;
mem_array[12619] = 16'hb9e1;
mem_array[12618] = 16'h3dc8;
mem_array[12621] = 16'h094d;
mem_array[12620] = 16'h3caa;
mem_array[12623] = 16'haaaf;
mem_array[12622] = 16'h3da9;
mem_array[12625] = 16'h6ccf;
mem_array[12624] = 16'hbe17;
mem_array[12627] = 16'h96b1;
mem_array[12626] = 16'h3e2e;
mem_array[12629] = 16'h9c44;
mem_array[12628] = 16'hbe57;
mem_array[12631] = 16'h8d3a;
mem_array[12630] = 16'hbe9c;
mem_array[12633] = 16'hc6d0;
mem_array[12632] = 16'hbd25;
mem_array[12635] = 16'h1a35;
mem_array[12634] = 16'hbf8e;
mem_array[12637] = 16'h74cf;
mem_array[12636] = 16'h3e1e;
mem_array[12639] = 16'headc;
mem_array[12638] = 16'hbe2a;
mem_array[12641] = 16'hf718;
mem_array[12640] = 16'hbe1d;
mem_array[12643] = 16'h51a6;
mem_array[12642] = 16'h3d6c;
mem_array[12645] = 16'h30b4;
mem_array[12644] = 16'hbddd;
mem_array[12647] = 16'hdfe8;
mem_array[12646] = 16'hbd19;
mem_array[12649] = 16'h3baf;
mem_array[12648] = 16'h3e71;
mem_array[12651] = 16'h5da3;
mem_array[12650] = 16'hbef5;
mem_array[12653] = 16'h981a;
mem_array[12652] = 16'h3c66;
mem_array[12655] = 16'h3996;
mem_array[12654] = 16'hbea1;
mem_array[12657] = 16'hd535;
mem_array[12656] = 16'hbd1a;
mem_array[12659] = 16'hcf13;
mem_array[12658] = 16'hbe9b;
mem_array[12661] = 16'h74bb;
mem_array[12660] = 16'hbe81;
mem_array[12663] = 16'h6b54;
mem_array[12662] = 16'hbe31;
mem_array[12665] = 16'h538c;
mem_array[12664] = 16'h3d2c;
mem_array[12667] = 16'h1c05;
mem_array[12666] = 16'h3dc0;
mem_array[12669] = 16'h15fd;
mem_array[12668] = 16'hbe9d;
mem_array[12671] = 16'h2463;
mem_array[12670] = 16'hbea0;
mem_array[12673] = 16'ha664;
mem_array[12672] = 16'hbedc;
mem_array[12675] = 16'h5a9a;
mem_array[12674] = 16'h3ded;
mem_array[12677] = 16'h2ed1;
mem_array[12676] = 16'hbe74;
mem_array[12679] = 16'h9e42;
mem_array[12678] = 16'h3d2d;
mem_array[12681] = 16'h01d4;
mem_array[12680] = 16'h3d3c;
mem_array[12683] = 16'h1894;
mem_array[12682] = 16'hbbbc;
mem_array[12685] = 16'h2a70;
mem_array[12684] = 16'hbe59;
mem_array[12687] = 16'h22f0;
mem_array[12686] = 16'h3e11;
mem_array[12689] = 16'h885a;
mem_array[12688] = 16'h3db5;
mem_array[12691] = 16'hfe51;
mem_array[12690] = 16'hbd0f;
mem_array[12693] = 16'h06c1;
mem_array[12692] = 16'hbee0;
mem_array[12695] = 16'hf601;
mem_array[12694] = 16'hbf90;
mem_array[12697] = 16'h6f6f;
mem_array[12696] = 16'h3c21;
mem_array[12699] = 16'hc4d5;
mem_array[12698] = 16'hbeb1;
mem_array[12701] = 16'ha0ac;
mem_array[12700] = 16'hbc8b;
mem_array[12703] = 16'hd27f;
mem_array[12702] = 16'h3ca1;
mem_array[12705] = 16'ha55f;
mem_array[12704] = 16'hbdf0;
mem_array[12707] = 16'h0b19;
mem_array[12706] = 16'hbd1a;
mem_array[12709] = 16'h1b60;
mem_array[12708] = 16'hbe01;
mem_array[12711] = 16'h1e88;
mem_array[12710] = 16'hbf0f;
mem_array[12713] = 16'h08f8;
mem_array[12712] = 16'h3d6f;
mem_array[12715] = 16'h2d9c;
mem_array[12714] = 16'hbefd;
mem_array[12717] = 16'h0029;
mem_array[12716] = 16'h3d78;
mem_array[12719] = 16'heef5;
mem_array[12718] = 16'hbf07;
mem_array[12721] = 16'h9c00;
mem_array[12720] = 16'h3d90;
mem_array[12723] = 16'h406e;
mem_array[12722] = 16'hbe33;
mem_array[12725] = 16'h7d79;
mem_array[12724] = 16'h3dde;
mem_array[12727] = 16'ha61e;
mem_array[12726] = 16'hbd02;
mem_array[12729] = 16'h516f;
mem_array[12728] = 16'hbe86;
mem_array[12731] = 16'h5c2b;
mem_array[12730] = 16'h3d61;
mem_array[12733] = 16'hef92;
mem_array[12732] = 16'h3d87;
mem_array[12735] = 16'h8db9;
mem_array[12734] = 16'hbbc1;
mem_array[12737] = 16'h6232;
mem_array[12736] = 16'hbee5;
mem_array[12739] = 16'hfc4a;
mem_array[12738] = 16'hbd33;
mem_array[12741] = 16'hcad8;
mem_array[12740] = 16'hbe09;
mem_array[12743] = 16'hda3f;
mem_array[12742] = 16'hbd8e;
mem_array[12745] = 16'h3d7d;
mem_array[12744] = 16'hbf26;
mem_array[12747] = 16'hbeec;
mem_array[12746] = 16'h3e2f;
mem_array[12749] = 16'hcdcc;
mem_array[12748] = 16'hbe0c;
mem_array[12751] = 16'hfb9d;
mem_array[12750] = 16'hbe1d;
mem_array[12753] = 16'hd340;
mem_array[12752] = 16'hbdb8;
mem_array[12755] = 16'h5bcc;
mem_array[12754] = 16'hbeea;
mem_array[12757] = 16'h260d;
mem_array[12756] = 16'h3e8f;
mem_array[12759] = 16'h6d69;
mem_array[12758] = 16'hbe9d;
mem_array[12761] = 16'h5e8a;
mem_array[12760] = 16'hbe09;
mem_array[12763] = 16'h5fd6;
mem_array[12762] = 16'hbdd9;
mem_array[12765] = 16'he131;
mem_array[12764] = 16'hbf16;
mem_array[12767] = 16'he64b;
mem_array[12766] = 16'hbe48;
mem_array[12769] = 16'hb273;
mem_array[12768] = 16'hbe00;
mem_array[12771] = 16'h8ef8;
mem_array[12770] = 16'hbe83;
mem_array[12773] = 16'h0429;
mem_array[12772] = 16'hbd1e;
mem_array[12775] = 16'h6729;
mem_array[12774] = 16'hbe43;
mem_array[12777] = 16'hd366;
mem_array[12776] = 16'h3e7a;
mem_array[12779] = 16'h91bf;
mem_array[12778] = 16'hbe23;
mem_array[12781] = 16'h78e0;
mem_array[12780] = 16'h3e13;
mem_array[12783] = 16'h8cb0;
mem_array[12782] = 16'hbe98;
mem_array[12785] = 16'h917b;
mem_array[12784] = 16'hbbeb;
mem_array[12787] = 16'h27ee;
mem_array[12786] = 16'h3ebf;
mem_array[12789] = 16'hb920;
mem_array[12788] = 16'hbeda;
mem_array[12791] = 16'h2845;
mem_array[12790] = 16'h3cdb;
mem_array[12793] = 16'ha3e1;
mem_array[12792] = 16'h3dbb;
mem_array[12795] = 16'h3e5f;
mem_array[12794] = 16'hbe28;
mem_array[12797] = 16'h60c3;
mem_array[12796] = 16'hbe1a;
mem_array[12799] = 16'h5192;
mem_array[12798] = 16'hbe7b;
mem_array[12801] = 16'h60f3;
mem_array[12800] = 16'hbbf6;
mem_array[12803] = 16'h29aa;
mem_array[12802] = 16'h3d28;
mem_array[12805] = 16'h18bd;
mem_array[12804] = 16'hbed0;
mem_array[12807] = 16'hcd11;
mem_array[12806] = 16'h3d60;
mem_array[12809] = 16'h3315;
mem_array[12808] = 16'hbe69;
mem_array[12811] = 16'hc0e4;
mem_array[12810] = 16'hbe82;
mem_array[12813] = 16'hd16c;
mem_array[12812] = 16'h3e6f;
mem_array[12815] = 16'h337e;
mem_array[12814] = 16'hbd5b;
mem_array[12817] = 16'h8b7a;
mem_array[12816] = 16'h3e8b;
mem_array[12819] = 16'hdba4;
mem_array[12818] = 16'hbe4f;
mem_array[12821] = 16'h786a;
mem_array[12820] = 16'hbe08;
mem_array[12823] = 16'heb24;
mem_array[12822] = 16'hbd09;
mem_array[12825] = 16'hff0e;
mem_array[12824] = 16'h3e60;
mem_array[12827] = 16'hfd19;
mem_array[12826] = 16'hbea4;
mem_array[12829] = 16'hb9b1;
mem_array[12828] = 16'h3e05;
mem_array[12831] = 16'h0bdf;
mem_array[12830] = 16'h3d80;
mem_array[12833] = 16'hccaa;
mem_array[12832] = 16'hbd0c;
mem_array[12835] = 16'hc626;
mem_array[12834] = 16'hbe8e;
mem_array[12837] = 16'h1eb7;
mem_array[12836] = 16'h3db6;
mem_array[12839] = 16'hedd7;
mem_array[12838] = 16'hbe1c;
mem_array[12841] = 16'h504f;
mem_array[12840] = 16'hbd71;
mem_array[12843] = 16'h47aa;
mem_array[12842] = 16'hbe55;
mem_array[12845] = 16'hf02e;
mem_array[12844] = 16'hbd33;
mem_array[12847] = 16'h7831;
mem_array[12846] = 16'h3f13;
mem_array[12849] = 16'h2716;
mem_array[12848] = 16'h3cdf;
mem_array[12851] = 16'h7112;
mem_array[12850] = 16'h3ed1;
mem_array[12853] = 16'hcc47;
mem_array[12852] = 16'hbe86;
mem_array[12855] = 16'h8fbc;
mem_array[12854] = 16'hbe36;
mem_array[12857] = 16'h578e;
mem_array[12856] = 16'hbe8b;
mem_array[12859] = 16'hbd71;
mem_array[12858] = 16'hbd0e;
mem_array[12861] = 16'h294d;
mem_array[12860] = 16'hbdb1;
mem_array[12863] = 16'h2180;
mem_array[12862] = 16'hbd1c;
mem_array[12865] = 16'h20c4;
mem_array[12864] = 16'hbe06;
mem_array[12867] = 16'hc2d7;
mem_array[12866] = 16'hbde0;
mem_array[12869] = 16'hbc5e;
mem_array[12868] = 16'h3df8;
mem_array[12871] = 16'h052c;
mem_array[12870] = 16'hbe14;
mem_array[12873] = 16'h7bec;
mem_array[12872] = 16'h3e30;
mem_array[12875] = 16'h4762;
mem_array[12874] = 16'h3e5b;
mem_array[12877] = 16'h251c;
mem_array[12876] = 16'hbdf3;
mem_array[12879] = 16'hf85a;
mem_array[12878] = 16'hbec4;
mem_array[12881] = 16'h118f;
mem_array[12880] = 16'hbed1;
mem_array[12883] = 16'hf5e0;
mem_array[12882] = 16'hbcff;
mem_array[12885] = 16'h2f1b;
mem_array[12884] = 16'hbdf6;
mem_array[12887] = 16'h7eae;
mem_array[12886] = 16'hbe11;
mem_array[12889] = 16'hb3b9;
mem_array[12888] = 16'h3d84;
mem_array[12891] = 16'hbfe3;
mem_array[12890] = 16'hbda8;
mem_array[12893] = 16'h16ad;
mem_array[12892] = 16'h3dfb;
mem_array[12895] = 16'hc30d;
mem_array[12894] = 16'hbdaf;
mem_array[12897] = 16'haeac;
mem_array[12896] = 16'hbe82;
mem_array[12899] = 16'he395;
mem_array[12898] = 16'hbefd;
mem_array[12901] = 16'h9b52;
mem_array[12900] = 16'h3e20;
mem_array[12903] = 16'haf05;
mem_array[12902] = 16'h3d78;
mem_array[12905] = 16'h5c34;
mem_array[12904] = 16'h3e38;
mem_array[12907] = 16'h4d8c;
mem_array[12906] = 16'h3eb1;
mem_array[12909] = 16'h1ba0;
mem_array[12908] = 16'h3ddd;
mem_array[12911] = 16'hc31c;
mem_array[12910] = 16'h3d6f;
mem_array[12913] = 16'h2ae6;
mem_array[12912] = 16'hbcdb;
mem_array[12915] = 16'hd417;
mem_array[12914] = 16'hbdae;
mem_array[12917] = 16'h3523;
mem_array[12916] = 16'hbc07;
mem_array[12919] = 16'hfc60;
mem_array[12918] = 16'hbe1e;
mem_array[12921] = 16'h06c2;
mem_array[12920] = 16'hbd8d;
mem_array[12923] = 16'h5689;
mem_array[12922] = 16'h3d13;
mem_array[12925] = 16'h7496;
mem_array[12924] = 16'hbde0;
mem_array[12927] = 16'hdfbb;
mem_array[12926] = 16'hbe92;
mem_array[12929] = 16'hc126;
mem_array[12928] = 16'h3ebe;
mem_array[12931] = 16'hbf1d;
mem_array[12930] = 16'h3baa;
mem_array[12933] = 16'h0420;
mem_array[12932] = 16'h3e3a;
mem_array[12935] = 16'h876e;
mem_array[12934] = 16'h3ea0;
mem_array[12937] = 16'ha451;
mem_array[12936] = 16'h3d66;
mem_array[12939] = 16'hf057;
mem_array[12938] = 16'hbd77;
mem_array[12941] = 16'he43e;
mem_array[12940] = 16'hbe93;
mem_array[12943] = 16'hd57c;
mem_array[12942] = 16'hbd59;
mem_array[12945] = 16'ha8f1;
mem_array[12944] = 16'hbee4;
mem_array[12947] = 16'hd3b7;
mem_array[12946] = 16'hbe14;
mem_array[12949] = 16'hfca9;
mem_array[12948] = 16'hbce8;
mem_array[12951] = 16'h57f5;
mem_array[12950] = 16'h3d17;
mem_array[12953] = 16'h9459;
mem_array[12952] = 16'hbda6;
mem_array[12955] = 16'h363a;
mem_array[12954] = 16'hbdb4;
mem_array[12957] = 16'h4049;
mem_array[12956] = 16'hbc13;
mem_array[12959] = 16'hdda9;
mem_array[12958] = 16'hbe91;
mem_array[12961] = 16'hb583;
mem_array[12960] = 16'hbe65;
mem_array[12963] = 16'h1638;
mem_array[12962] = 16'hbe46;
mem_array[12965] = 16'hbaaf;
mem_array[12964] = 16'hbe80;
mem_array[12967] = 16'hfb6b;
mem_array[12966] = 16'hbe1d;
mem_array[12969] = 16'h98e5;
mem_array[12968] = 16'h3e17;
mem_array[12971] = 16'haf5a;
mem_array[12970] = 16'h3dee;
mem_array[12973] = 16'hdbd0;
mem_array[12972] = 16'hbe85;
mem_array[12975] = 16'h1138;
mem_array[12974] = 16'hbd4d;
mem_array[12977] = 16'hc308;
mem_array[12976] = 16'h3cd9;
mem_array[12979] = 16'he808;
mem_array[12978] = 16'hbf68;
mem_array[12981] = 16'h7af7;
mem_array[12980] = 16'h3b80;
mem_array[12983] = 16'h85ec;
mem_array[12982] = 16'h3d89;
mem_array[12985] = 16'h9f80;
mem_array[12984] = 16'hbd2d;
mem_array[12987] = 16'hc6f0;
mem_array[12986] = 16'hbead;
mem_array[12989] = 16'hd260;
mem_array[12988] = 16'h3dd5;
mem_array[12991] = 16'h148e;
mem_array[12990] = 16'h3e3a;
mem_array[12993] = 16'h4916;
mem_array[12992] = 16'h3b88;
mem_array[12995] = 16'hc06e;
mem_array[12994] = 16'h3ce0;
mem_array[12997] = 16'h13f4;
mem_array[12996] = 16'h3e5e;
mem_array[12999] = 16'h4e64;
mem_array[12998] = 16'h3e98;
mem_array[13001] = 16'h923e;
mem_array[13000] = 16'h3e27;
mem_array[13003] = 16'hde0a;
mem_array[13002] = 16'hbdb5;
mem_array[13005] = 16'h07dd;
mem_array[13004] = 16'hbf1d;
mem_array[13007] = 16'h8776;
mem_array[13006] = 16'hbe9b;
mem_array[13009] = 16'hdeb5;
mem_array[13008] = 16'h3d99;
mem_array[13011] = 16'h1f3f;
mem_array[13010] = 16'hbea8;
mem_array[13013] = 16'h878b;
mem_array[13012] = 16'hbe1b;
mem_array[13015] = 16'h3fec;
mem_array[13014] = 16'h3e9c;
mem_array[13017] = 16'hdb55;
mem_array[13016] = 16'h3dad;
mem_array[13019] = 16'h0640;
mem_array[13018] = 16'hbc9b;
mem_array[13021] = 16'h2752;
mem_array[13020] = 16'h3e4e;
mem_array[13023] = 16'h64c6;
mem_array[13022] = 16'hbeb7;
mem_array[13025] = 16'he139;
mem_array[13024] = 16'hbea4;
mem_array[13027] = 16'h7220;
mem_array[13026] = 16'hbeef;
mem_array[13029] = 16'hecee;
mem_array[13028] = 16'hbcb2;
mem_array[13031] = 16'h0e9b;
mem_array[13030] = 16'h3e3b;
mem_array[13033] = 16'hd3d5;
mem_array[13032] = 16'hbe3d;
mem_array[13035] = 16'h461e;
mem_array[13034] = 16'hbe60;
mem_array[13037] = 16'h3671;
mem_array[13036] = 16'hbe58;
mem_array[13039] = 16'h908a;
mem_array[13038] = 16'hbec8;
mem_array[13041] = 16'h6145;
mem_array[13040] = 16'hbd95;
mem_array[13043] = 16'h000c;
mem_array[13042] = 16'h3d89;
mem_array[13045] = 16'h63d3;
mem_array[13044] = 16'hbe59;
mem_array[13047] = 16'hb9fe;
mem_array[13046] = 16'hbe7d;
mem_array[13049] = 16'ha58a;
mem_array[13048] = 16'h3ecd;
mem_array[13051] = 16'h5455;
mem_array[13050] = 16'h3e22;
mem_array[13053] = 16'h7c2f;
mem_array[13052] = 16'h3dce;
mem_array[13055] = 16'h83e9;
mem_array[13054] = 16'hbe00;
mem_array[13057] = 16'h0fce;
mem_array[13056] = 16'hbe07;
mem_array[13059] = 16'h59aa;
mem_array[13058] = 16'h3da2;
mem_array[13061] = 16'h8a2d;
mem_array[13060] = 16'h3d53;
mem_array[13063] = 16'h64b3;
mem_array[13062] = 16'h3e5f;
mem_array[13065] = 16'hebd8;
mem_array[13064] = 16'hbeb0;
mem_array[13067] = 16'h6ad3;
mem_array[13066] = 16'hbeab;
mem_array[13069] = 16'h0d4a;
mem_array[13068] = 16'hbe96;
mem_array[13071] = 16'hb9a4;
mem_array[13070] = 16'hbe37;
mem_array[13073] = 16'h66fd;
mem_array[13072] = 16'hbc42;
mem_array[13075] = 16'h16e4;
mem_array[13074] = 16'h3eb1;
mem_array[13077] = 16'hb492;
mem_array[13076] = 16'h3d87;
mem_array[13079] = 16'hd22f;
mem_array[13078] = 16'h3e8d;
mem_array[13081] = 16'hc3f1;
mem_array[13080] = 16'hbe42;
mem_array[13083] = 16'h6870;
mem_array[13082] = 16'hbf00;
mem_array[13085] = 16'h89e9;
mem_array[13084] = 16'h3e09;
mem_array[13087] = 16'h4b03;
mem_array[13086] = 16'hbd97;
mem_array[13089] = 16'h0eb4;
mem_array[13088] = 16'hbdf1;
mem_array[13091] = 16'h5c46;
mem_array[13090] = 16'h3e98;
mem_array[13093] = 16'h5a58;
mem_array[13092] = 16'hbea1;
mem_array[13095] = 16'hdb19;
mem_array[13094] = 16'h3e39;
mem_array[13097] = 16'h39c2;
mem_array[13096] = 16'h3e9f;
mem_array[13099] = 16'h6774;
mem_array[13098] = 16'hbee8;
mem_array[13101] = 16'h3140;
mem_array[13100] = 16'h3c96;
mem_array[13103] = 16'hafb3;
mem_array[13102] = 16'hbd59;
mem_array[13105] = 16'h0ca8;
mem_array[13104] = 16'hbe51;
mem_array[13107] = 16'h5aee;
mem_array[13106] = 16'h3ec3;
mem_array[13109] = 16'h074c;
mem_array[13108] = 16'h3ebd;
mem_array[13111] = 16'h4887;
mem_array[13110] = 16'hbca2;
mem_array[13113] = 16'h8a5c;
mem_array[13112] = 16'h3e27;
mem_array[13115] = 16'haafe;
mem_array[13114] = 16'h3ec7;
mem_array[13117] = 16'h9e6b;
mem_array[13116] = 16'hbccb;
mem_array[13119] = 16'h2435;
mem_array[13118] = 16'h3ed0;
mem_array[13121] = 16'hf17b;
mem_array[13120] = 16'h3d8a;
mem_array[13123] = 16'hced1;
mem_array[13122] = 16'h3da8;
mem_array[13125] = 16'h3d18;
mem_array[13124] = 16'hbf4a;
mem_array[13127] = 16'h287b;
mem_array[13126] = 16'hbec1;
mem_array[13129] = 16'hf4b2;
mem_array[13128] = 16'h3d82;
mem_array[13131] = 16'h6257;
mem_array[13130] = 16'h3d61;
mem_array[13133] = 16'h9baf;
mem_array[13132] = 16'h3e81;
mem_array[13135] = 16'h5cb4;
mem_array[13134] = 16'h3ef6;
mem_array[13137] = 16'haa01;
mem_array[13136] = 16'h3efd;
mem_array[13139] = 16'h12ee;
mem_array[13138] = 16'h3eaa;
mem_array[13141] = 16'hf18a;
mem_array[13140] = 16'hbe00;
mem_array[13143] = 16'he299;
mem_array[13142] = 16'hbc9c;
mem_array[13145] = 16'hd623;
mem_array[13144] = 16'hbf22;
mem_array[13147] = 16'hfb61;
mem_array[13146] = 16'h3da9;
mem_array[13149] = 16'h06fa;
mem_array[13148] = 16'h3f02;
mem_array[13151] = 16'h52a1;
mem_array[13150] = 16'h3ea3;
mem_array[13153] = 16'h1cd9;
mem_array[13152] = 16'hbf76;
mem_array[13155] = 16'hf642;
mem_array[13154] = 16'h3e14;
mem_array[13157] = 16'h56f6;
mem_array[13156] = 16'hbf20;
mem_array[13159] = 16'hb1b5;
mem_array[13158] = 16'hbf87;
mem_array[13161] = 16'hf0ad;
mem_array[13160] = 16'h3d41;
mem_array[13163] = 16'h35f0;
mem_array[13162] = 16'hbc67;
mem_array[13165] = 16'h6646;
mem_array[13164] = 16'hbf1c;
mem_array[13167] = 16'h9908;
mem_array[13166] = 16'hbd92;
mem_array[13169] = 16'hf247;
mem_array[13168] = 16'hbe02;
mem_array[13171] = 16'h671a;
mem_array[13170] = 16'h3e1a;
mem_array[13173] = 16'heade;
mem_array[13172] = 16'hbeea;
mem_array[13175] = 16'h8d4d;
mem_array[13174] = 16'h3ea2;
mem_array[13177] = 16'h4576;
mem_array[13176] = 16'hbf0d;
mem_array[13179] = 16'hb6d8;
mem_array[13178] = 16'h3ea3;
mem_array[13181] = 16'h9cac;
mem_array[13180] = 16'h3ef7;
mem_array[13183] = 16'h2e41;
mem_array[13182] = 16'hbe83;
mem_array[13185] = 16'h98c1;
mem_array[13184] = 16'hbf19;
mem_array[13187] = 16'hb74d;
mem_array[13186] = 16'hbeb6;
mem_array[13189] = 16'h0da6;
mem_array[13188] = 16'hbee9;
mem_array[13191] = 16'h756e;
mem_array[13190] = 16'h3ea6;
mem_array[13193] = 16'hb109;
mem_array[13192] = 16'h3e55;
mem_array[13195] = 16'h39b8;
mem_array[13194] = 16'h3edd;
mem_array[13197] = 16'h05a9;
mem_array[13196] = 16'hbf44;
mem_array[13199] = 16'hb680;
mem_array[13198] = 16'h3d5d;
mem_array[13201] = 16'h0daa;
mem_array[13200] = 16'hbfd0;
mem_array[13203] = 16'hd7d7;
mem_array[13202] = 16'hbea1;
mem_array[13205] = 16'hf081;
mem_array[13204] = 16'hbf1f;
mem_array[13207] = 16'h1c10;
mem_array[13206] = 16'hbf28;
mem_array[13209] = 16'h9f7d;
mem_array[13208] = 16'h3df8;
mem_array[13211] = 16'h96f0;
mem_array[13210] = 16'h3f04;
mem_array[13213] = 16'h4309;
mem_array[13212] = 16'hc00c;
mem_array[13215] = 16'h8ab4;
mem_array[13214] = 16'h3df3;
mem_array[13217] = 16'h183a;
mem_array[13216] = 16'hbfb9;
mem_array[13219] = 16'h32bd;
mem_array[13218] = 16'hbf5b;
mem_array[13221] = 16'hfb65;
mem_array[13220] = 16'hbd96;
mem_array[13223] = 16'hfd5a;
mem_array[13222] = 16'h38f3;
mem_array[13225] = 16'h31f0;
mem_array[13224] = 16'hbf38;
mem_array[13227] = 16'hfede;
mem_array[13226] = 16'hbe5a;
mem_array[13229] = 16'h0b70;
mem_array[13228] = 16'hbf05;
mem_array[13231] = 16'hc020;
mem_array[13230] = 16'hbee2;
mem_array[13233] = 16'hec51;
mem_array[13232] = 16'hbf31;
mem_array[13235] = 16'h7d2e;
mem_array[13234] = 16'hbeca;
mem_array[13237] = 16'h0fdc;
mem_array[13236] = 16'hbf58;
mem_array[13239] = 16'h5913;
mem_array[13238] = 16'hbe5c;
mem_array[13241] = 16'h60aa;
mem_array[13240] = 16'h3ea4;
mem_array[13243] = 16'h02b0;
mem_array[13242] = 16'hbc2b;
mem_array[13245] = 16'hbb82;
mem_array[13244] = 16'hbf99;
mem_array[13247] = 16'hf26d;
mem_array[13246] = 16'hbe58;
mem_array[13249] = 16'h4735;
mem_array[13248] = 16'hbeb5;
mem_array[13251] = 16'h26de;
mem_array[13250] = 16'h3eb4;
mem_array[13253] = 16'h4972;
mem_array[13252] = 16'h3f2c;
mem_array[13255] = 16'h811f;
mem_array[13254] = 16'h3e2a;
mem_array[13257] = 16'h4444;
mem_array[13256] = 16'hbf62;
mem_array[13259] = 16'h57e3;
mem_array[13258] = 16'hbf46;
mem_array[13261] = 16'hb8e1;
mem_array[13260] = 16'hc006;
mem_array[13263] = 16'h280d;
mem_array[13262] = 16'hbf0e;
mem_array[13265] = 16'hf4ee;
mem_array[13264] = 16'hbf85;
mem_array[13267] = 16'h91f2;
mem_array[13266] = 16'hbff3;
mem_array[13269] = 16'ha7e3;
mem_array[13268] = 16'hbdd9;
mem_array[13271] = 16'h2315;
mem_array[13270] = 16'h3f07;
mem_array[13273] = 16'ha710;
mem_array[13272] = 16'hbfae;
mem_array[13275] = 16'hb1df;
mem_array[13274] = 16'hbe91;
mem_array[13277] = 16'h1f7e;
mem_array[13276] = 16'hbeeb;
mem_array[13279] = 16'h4ba2;
mem_array[13278] = 16'hbeb6;
mem_array[13281] = 16'h2ae6;
mem_array[13280] = 16'h3cda;
mem_array[13283] = 16'h5596;
mem_array[13282] = 16'hbd04;
mem_array[13285] = 16'hbeb8;
mem_array[13284] = 16'hbef3;
mem_array[13287] = 16'h245f;
mem_array[13286] = 16'hbecb;
mem_array[13289] = 16'h92fb;
mem_array[13288] = 16'hbfb0;
mem_array[13291] = 16'h8aa5;
mem_array[13290] = 16'hbedb;
mem_array[13293] = 16'h03a0;
mem_array[13292] = 16'hbf8c;
mem_array[13295] = 16'h68a4;
mem_array[13294] = 16'hbeb4;
mem_array[13297] = 16'h84f8;
mem_array[13296] = 16'hbf0f;
mem_array[13299] = 16'hfe11;
mem_array[13298] = 16'hbe82;
mem_array[13301] = 16'h20f9;
mem_array[13300] = 16'hbe58;
mem_array[13303] = 16'ha2a9;
mem_array[13302] = 16'h3e22;
mem_array[13305] = 16'h105a;
mem_array[13304] = 16'hbebb;
mem_array[13307] = 16'h8244;
mem_array[13306] = 16'hbda2;
mem_array[13309] = 16'h484b;
mem_array[13308] = 16'hbf98;
mem_array[13311] = 16'he876;
mem_array[13310] = 16'hbf8f;
mem_array[13313] = 16'h7545;
mem_array[13312] = 16'h3f4c;
mem_array[13315] = 16'h195d;
mem_array[13314] = 16'h3d0f;
mem_array[13317] = 16'he265;
mem_array[13316] = 16'hbef5;
mem_array[13319] = 16'hc58e;
mem_array[13318] = 16'hbfb2;
mem_array[13321] = 16'h7180;
mem_array[13320] = 16'hbf4e;
mem_array[13323] = 16'hc9bd;
mem_array[13322] = 16'hbf13;
mem_array[13325] = 16'h6af9;
mem_array[13324] = 16'h3e2e;
mem_array[13327] = 16'h4969;
mem_array[13326] = 16'hbfe1;
mem_array[13329] = 16'h76fe;
mem_array[13328] = 16'h3eba;
mem_array[13331] = 16'h79bd;
mem_array[13330] = 16'h3e57;
mem_array[13333] = 16'hfd35;
mem_array[13332] = 16'hbe91;
mem_array[13335] = 16'h4f21;
mem_array[13334] = 16'h3eb9;
mem_array[13337] = 16'h4f88;
mem_array[13336] = 16'h3c1b;
mem_array[13339] = 16'h1acc;
mem_array[13338] = 16'h3e48;
mem_array[13341] = 16'h1d52;
mem_array[13340] = 16'hbcf5;
mem_array[13343] = 16'hc0fb;
mem_array[13342] = 16'h3d20;
mem_array[13345] = 16'h3641;
mem_array[13344] = 16'h3eeb;
mem_array[13347] = 16'h360c;
mem_array[13346] = 16'h3e10;
mem_array[13349] = 16'h3bcc;
mem_array[13348] = 16'hbeaa;
mem_array[13351] = 16'h45e7;
mem_array[13350] = 16'h3e4e;
mem_array[13353] = 16'h60a3;
mem_array[13352] = 16'h3dbb;
mem_array[13355] = 16'h406a;
mem_array[13354] = 16'hbe5e;
mem_array[13357] = 16'h9642;
mem_array[13356] = 16'hbeeb;
mem_array[13359] = 16'heb34;
mem_array[13358] = 16'h3e93;
mem_array[13361] = 16'h2982;
mem_array[13360] = 16'h3f3b;
mem_array[13363] = 16'h425e;
mem_array[13362] = 16'hbe3a;
mem_array[13365] = 16'h9381;
mem_array[13364] = 16'hbf09;
mem_array[13367] = 16'hed03;
mem_array[13366] = 16'hbf00;
mem_array[13369] = 16'h738f;
mem_array[13368] = 16'hbedf;
mem_array[13371] = 16'he4ca;
mem_array[13370] = 16'hbea6;
mem_array[13373] = 16'h35a4;
mem_array[13372] = 16'hbd73;
mem_array[13375] = 16'hde4f;
mem_array[13374] = 16'h3f31;
mem_array[13377] = 16'heac3;
mem_array[13376] = 16'h3bd8;
mem_array[13379] = 16'h2569;
mem_array[13378] = 16'hbfa6;
mem_array[13381] = 16'h3e61;
mem_array[13380] = 16'h3e62;
mem_array[13383] = 16'ha202;
mem_array[13382] = 16'hbf28;
mem_array[13385] = 16'h25f2;
mem_array[13384] = 16'h3dd8;
mem_array[13387] = 16'h3918;
mem_array[13386] = 16'hbf2e;
mem_array[13389] = 16'hcf2d;
mem_array[13388] = 16'hbf16;
mem_array[13391] = 16'h7d99;
mem_array[13390] = 16'h3f35;
mem_array[13393] = 16'h8aeb;
mem_array[13392] = 16'h3df4;
mem_array[13395] = 16'h1d83;
mem_array[13394] = 16'h3ea7;
mem_array[13397] = 16'hcada;
mem_array[13396] = 16'hbda8;
mem_array[13399] = 16'h4c98;
mem_array[13398] = 16'h3e92;
mem_array[13401] = 16'h8329;
mem_array[13400] = 16'h3d9b;
mem_array[13403] = 16'h09a7;
mem_array[13402] = 16'hbd3a;
mem_array[13405] = 16'hea07;
mem_array[13404] = 16'hbeb0;
mem_array[13407] = 16'h8e30;
mem_array[13406] = 16'hbd99;
mem_array[13409] = 16'h142d;
mem_array[13408] = 16'hbdc2;
mem_array[13411] = 16'h269c;
mem_array[13410] = 16'h3ef6;
mem_array[13413] = 16'h4d9f;
mem_array[13412] = 16'h3d4c;
mem_array[13415] = 16'h50f1;
mem_array[13414] = 16'h3e1d;
mem_array[13417] = 16'h67dd;
mem_array[13416] = 16'hbe58;
mem_array[13419] = 16'h0a06;
mem_array[13418] = 16'hbe9c;
mem_array[13421] = 16'h1e55;
mem_array[13420] = 16'hbf39;
mem_array[13423] = 16'hca48;
mem_array[13422] = 16'h3f63;
mem_array[13425] = 16'h4ae1;
mem_array[13424] = 16'hbc49;
mem_array[13427] = 16'h6bc6;
mem_array[13426] = 16'hbfc5;
mem_array[13429] = 16'hc57a;
mem_array[13428] = 16'hbe2a;
mem_array[13431] = 16'h2f86;
mem_array[13430] = 16'hbd3e;
mem_array[13433] = 16'h2ec0;
mem_array[13432] = 16'h3edf;
mem_array[13435] = 16'h8e7e;
mem_array[13434] = 16'h3fba;
mem_array[13437] = 16'h7234;
mem_array[13436] = 16'h3dca;
mem_array[13439] = 16'h60d8;
mem_array[13438] = 16'hbf47;
mem_array[13441] = 16'h8499;
mem_array[13440] = 16'h3da6;
mem_array[13443] = 16'h89bf;
mem_array[13442] = 16'h3f0c;
mem_array[13445] = 16'hbeea;
mem_array[13444] = 16'h3ea2;
mem_array[13447] = 16'hae51;
mem_array[13446] = 16'h3e5e;
mem_array[13449] = 16'hde75;
mem_array[13448] = 16'hbcc7;
mem_array[13451] = 16'he49d;
mem_array[13450] = 16'h3d9d;
mem_array[13453] = 16'h3e81;
mem_array[13452] = 16'hbc07;
mem_array[13455] = 16'hde1b;
mem_array[13454] = 16'h3e1c;
mem_array[13457] = 16'h1284;
mem_array[13456] = 16'hbbcb;
mem_array[13459] = 16'h86a8;
mem_array[13458] = 16'h3d46;
mem_array[13461] = 16'h4ce0;
mem_array[13460] = 16'h3cb3;
mem_array[13463] = 16'he280;
mem_array[13462] = 16'hbd44;
mem_array[13465] = 16'h4353;
mem_array[13464] = 16'h3ee7;
mem_array[13467] = 16'ha8d2;
mem_array[13466] = 16'hbd85;
mem_array[13469] = 16'ha9b0;
mem_array[13468] = 16'hbcda;
mem_array[13471] = 16'hb33a;
mem_array[13470] = 16'hbee3;
mem_array[13473] = 16'hdd03;
mem_array[13472] = 16'h3d48;
mem_array[13475] = 16'h6515;
mem_array[13474] = 16'h3d64;
mem_array[13477] = 16'h791c;
mem_array[13476] = 16'h3d0d;
mem_array[13479] = 16'h3bd7;
mem_array[13478] = 16'h3e0b;
mem_array[13481] = 16'h4b50;
mem_array[13480] = 16'hbd93;
mem_array[13483] = 16'haf5e;
mem_array[13482] = 16'h3dc8;
mem_array[13485] = 16'h2346;
mem_array[13484] = 16'hbddc;
mem_array[13487] = 16'hf0f4;
mem_array[13486] = 16'h3da9;
mem_array[13489] = 16'h24a9;
mem_array[13488] = 16'hbe0c;
mem_array[13491] = 16'hf2e7;
mem_array[13490] = 16'h3db6;
mem_array[13493] = 16'h6d85;
mem_array[13492] = 16'hbe85;
mem_array[13495] = 16'h8046;
mem_array[13494] = 16'h3c6f;
mem_array[13497] = 16'h660c;
mem_array[13496] = 16'hbc11;
mem_array[13499] = 16'h1875;
mem_array[13498] = 16'h3e42;
mem_array[13501] = 16'h26ad;
mem_array[13500] = 16'hbdde;
mem_array[13503] = 16'h68cf;
mem_array[13502] = 16'h3fb8;
mem_array[13505] = 16'h92f8;
mem_array[13504] = 16'h3f8f;
mem_array[13507] = 16'h4f07;
mem_array[13506] = 16'h3d1a;
mem_array[13509] = 16'h9c81;
mem_array[13508] = 16'h3f5e;
mem_array[13511] = 16'h1aa1;
mem_array[13510] = 16'h3df2;
mem_array[13513] = 16'h1e1d;
mem_array[13512] = 16'h3f27;
mem_array[13515] = 16'h3684;
mem_array[13514] = 16'h3f9f;
mem_array[13517] = 16'hab86;
mem_array[13516] = 16'h3fba;
mem_array[13519] = 16'hee40;
mem_array[13518] = 16'hbc83;
mem_array[13521] = 16'h98d4;
mem_array[13520] = 16'h3d31;
mem_array[13523] = 16'h302e;
mem_array[13522] = 16'hbc01;
mem_array[13525] = 16'h23ca;
mem_array[13524] = 16'hbf33;
mem_array[13527] = 16'h5145;
mem_array[13526] = 16'h3eab;
mem_array[13529] = 16'h9122;
mem_array[13528] = 16'h3f36;
mem_array[13531] = 16'hac38;
mem_array[13530] = 16'hbde8;
mem_array[13533] = 16'h3e85;
mem_array[13532] = 16'h3c96;
mem_array[13535] = 16'hc4e5;
mem_array[13534] = 16'hbe84;
mem_array[13537] = 16'h6082;
mem_array[13536] = 16'h3f66;
mem_array[13539] = 16'hdfc1;
mem_array[13538] = 16'h3e8f;
mem_array[13541] = 16'hce48;
mem_array[13540] = 16'hbf97;
mem_array[13543] = 16'hf159;
mem_array[13542] = 16'h3ea6;
mem_array[13545] = 16'h0577;
mem_array[13544] = 16'hbde4;
mem_array[13547] = 16'hd802;
mem_array[13546] = 16'hc004;
mem_array[13549] = 16'h6266;
mem_array[13548] = 16'hbee6;
mem_array[13551] = 16'hecee;
mem_array[13550] = 16'h4012;
mem_array[13553] = 16'haa5c;
mem_array[13552] = 16'hbda9;
mem_array[13555] = 16'h3320;
mem_array[13554] = 16'h3f4e;
mem_array[13557] = 16'hd0f7;
mem_array[13556] = 16'hbd44;
mem_array[13559] = 16'h9094;
mem_array[13558] = 16'hbfdf;
mem_array[13561] = 16'h84d1;
mem_array[13560] = 16'h3dce;
mem_array[13563] = 16'hd7fe;
mem_array[13562] = 16'h3f1a;
mem_array[13565] = 16'h89af;
mem_array[13564] = 16'hbcfd;
mem_array[13567] = 16'he27a;
mem_array[13566] = 16'h3e76;
mem_array[13569] = 16'h4a60;
mem_array[13568] = 16'h3e86;
mem_array[13571] = 16'hb1cc;
mem_array[13570] = 16'h3dd8;
mem_array[13573] = 16'he63e;
mem_array[13572] = 16'hbf63;
mem_array[13575] = 16'hcec5;
mem_array[13574] = 16'hbf3c;
mem_array[13577] = 16'hca8a;
mem_array[13576] = 16'hbe81;
mem_array[13579] = 16'h5570;
mem_array[13578] = 16'h3ef5;
mem_array[13581] = 16'h5636;
mem_array[13580] = 16'h3d2e;
mem_array[13583] = 16'h3ef1;
mem_array[13582] = 16'h3dc2;
mem_array[13585] = 16'h6bfd;
mem_array[13584] = 16'h3e90;
mem_array[13587] = 16'ha42e;
mem_array[13586] = 16'hbf96;
mem_array[13589] = 16'h2eec;
mem_array[13588] = 16'h3e9f;
mem_array[13591] = 16'h4fcf;
mem_array[13590] = 16'hbf32;
mem_array[13593] = 16'h5740;
mem_array[13592] = 16'hbdbd;
mem_array[13595] = 16'h95e2;
mem_array[13594] = 16'h3e8b;
mem_array[13597] = 16'hb946;
mem_array[13596] = 16'h3f7f;
mem_array[13599] = 16'h7c3d;
mem_array[13598] = 16'h3f09;
mem_array[13601] = 16'h945c;
mem_array[13600] = 16'h3ea0;
mem_array[13603] = 16'h92dc;
mem_array[13602] = 16'h3c38;
mem_array[13605] = 16'h4dc6;
mem_array[13604] = 16'hbbaa;
mem_array[13607] = 16'h441c;
mem_array[13606] = 16'hbec8;
mem_array[13609] = 16'hbe08;
mem_array[13608] = 16'hbdea;
mem_array[13611] = 16'h8c4f;
mem_array[13610] = 16'h3fd1;
mem_array[13613] = 16'hdc65;
mem_array[13612] = 16'hbef3;
mem_array[13615] = 16'hd1d6;
mem_array[13614] = 16'hbcc8;
mem_array[13617] = 16'h274c;
mem_array[13616] = 16'hbe26;
mem_array[13619] = 16'hdde1;
mem_array[13618] = 16'h3e0c;
mem_array[13621] = 16'h02ae;
mem_array[13620] = 16'h3f86;
mem_array[13623] = 16'hd43e;
mem_array[13622] = 16'h3f10;
mem_array[13625] = 16'h3d68;
mem_array[13624] = 16'h3f02;
mem_array[13627] = 16'hc3ed;
mem_array[13626] = 16'hbdd4;
mem_array[13629] = 16'h5262;
mem_array[13628] = 16'h3f4d;
mem_array[13631] = 16'hd27b;
mem_array[13630] = 16'hbdb0;
mem_array[13633] = 16'hf13a;
mem_array[13632] = 16'h3d34;
mem_array[13635] = 16'hd10b;
mem_array[13634] = 16'h3ead;
mem_array[13637] = 16'h368e;
mem_array[13636] = 16'hbf6f;
mem_array[13639] = 16'hc6ba;
mem_array[13638] = 16'h3ebf;
mem_array[13641] = 16'h719b;
mem_array[13640] = 16'h3d06;
mem_array[13643] = 16'hea55;
mem_array[13642] = 16'h3d21;
mem_array[13645] = 16'hfacf;
mem_array[13644] = 16'h3ed9;
mem_array[13647] = 16'h8ae8;
mem_array[13646] = 16'hbf92;
mem_array[13649] = 16'h9b6a;
mem_array[13648] = 16'hbde1;
mem_array[13651] = 16'h69ae;
mem_array[13650] = 16'hbe4d;
mem_array[13653] = 16'h3798;
mem_array[13652] = 16'hbf30;
mem_array[13655] = 16'hfa4f;
mem_array[13654] = 16'h3f06;
mem_array[13657] = 16'hef39;
mem_array[13656] = 16'h3e96;
mem_array[13659] = 16'h9d60;
mem_array[13658] = 16'h3e29;
mem_array[13661] = 16'hae75;
mem_array[13660] = 16'hbd6a;
mem_array[13663] = 16'h05cd;
mem_array[13662] = 16'h3e9b;
mem_array[13665] = 16'h7bb9;
mem_array[13664] = 16'hbf35;
mem_array[13667] = 16'h8ae6;
mem_array[13666] = 16'hbed5;
mem_array[13669] = 16'h5fec;
mem_array[13668] = 16'h3e0c;
mem_array[13671] = 16'h2423;
mem_array[13670] = 16'h3f63;
mem_array[13673] = 16'h816a;
mem_array[13672] = 16'h3e65;
mem_array[13675] = 16'h69ab;
mem_array[13674] = 16'hbd20;
mem_array[13677] = 16'hcd8f;
mem_array[13676] = 16'hbe42;
mem_array[13679] = 16'h1115;
mem_array[13678] = 16'hbf1c;
mem_array[13681] = 16'hb75a;
mem_array[13680] = 16'h3f2d;
mem_array[13683] = 16'h928d;
mem_array[13682] = 16'hbca7;
mem_array[13685] = 16'hafcc;
mem_array[13684] = 16'h3f07;
mem_array[13687] = 16'h5477;
mem_array[13686] = 16'hbd67;
mem_array[13689] = 16'h8aed;
mem_array[13688] = 16'hbf15;
mem_array[13691] = 16'h2342;
mem_array[13690] = 16'hbf2f;
mem_array[13693] = 16'had06;
mem_array[13692] = 16'h3f68;
mem_array[13695] = 16'hba97;
mem_array[13694] = 16'hbe17;
mem_array[13697] = 16'h29fb;
mem_array[13696] = 16'hbeee;
mem_array[13699] = 16'hca7d;
mem_array[13698] = 16'hbe1b;
mem_array[13701] = 16'hfa8e;
mem_array[13700] = 16'hbda1;
mem_array[13703] = 16'h8a29;
mem_array[13702] = 16'hbc6c;
mem_array[13705] = 16'h21e9;
mem_array[13704] = 16'hbee9;
mem_array[13707] = 16'hb33b;
mem_array[13706] = 16'hbe3f;
mem_array[13709] = 16'haa24;
mem_array[13708] = 16'h3e8b;
mem_array[13711] = 16'h2505;
mem_array[13710] = 16'h3e10;
mem_array[13713] = 16'h5159;
mem_array[13712] = 16'hbd15;
mem_array[13715] = 16'h14b1;
mem_array[13714] = 16'h3f01;
mem_array[13717] = 16'h8470;
mem_array[13716] = 16'hbe91;
mem_array[13719] = 16'h5510;
mem_array[13718] = 16'h3c6d;
mem_array[13721] = 16'h6550;
mem_array[13720] = 16'hbe14;
mem_array[13723] = 16'he49b;
mem_array[13722] = 16'hbe13;
mem_array[13725] = 16'hc869;
mem_array[13724] = 16'hbf69;
mem_array[13727] = 16'h4904;
mem_array[13726] = 16'hbdb7;
mem_array[13729] = 16'hdf3f;
mem_array[13728] = 16'h3dfa;
mem_array[13731] = 16'hcf24;
mem_array[13730] = 16'h3d3c;
mem_array[13733] = 16'h13b0;
mem_array[13732] = 16'h3bb8;
mem_array[13735] = 16'h00f0;
mem_array[13734] = 16'h3cc7;
mem_array[13737] = 16'hcd85;
mem_array[13736] = 16'hbec6;
mem_array[13739] = 16'h5d1d;
mem_array[13738] = 16'hbf07;
mem_array[13741] = 16'h9bae;
mem_array[13740] = 16'hbdd6;
mem_array[13743] = 16'h2bad;
mem_array[13742] = 16'hbc39;
mem_array[13745] = 16'h0612;
mem_array[13744] = 16'hbe4a;
mem_array[13747] = 16'h862e;
mem_array[13746] = 16'h3d1f;
mem_array[13749] = 16'h8876;
mem_array[13748] = 16'hbf8a;
mem_array[13751] = 16'h48e1;
mem_array[13750] = 16'hbea1;
mem_array[13753] = 16'ha08d;
mem_array[13752] = 16'h3e4f;
mem_array[13755] = 16'h42ca;
mem_array[13754] = 16'hbeb6;
mem_array[13757] = 16'hfe0a;
mem_array[13756] = 16'hbf01;
mem_array[13759] = 16'h449f;
mem_array[13758] = 16'hbba3;
mem_array[13761] = 16'h31c8;
mem_array[13760] = 16'h3bcd;
mem_array[13763] = 16'h9ecb;
mem_array[13762] = 16'hbcaf;
mem_array[13765] = 16'hd42b;
mem_array[13764] = 16'hbe5b;
mem_array[13767] = 16'hd5ca;
mem_array[13766] = 16'hbda3;
mem_array[13769] = 16'h5ee0;
mem_array[13768] = 16'hbdd4;
mem_array[13771] = 16'h413e;
mem_array[13770] = 16'h3e2f;
mem_array[13773] = 16'h3bc2;
mem_array[13772] = 16'h3dab;
mem_array[13775] = 16'hbbb4;
mem_array[13774] = 16'h3ea9;
mem_array[13777] = 16'hcd48;
mem_array[13776] = 16'hbd72;
mem_array[13779] = 16'haa67;
mem_array[13778] = 16'h3d25;
mem_array[13781] = 16'h3181;
mem_array[13780] = 16'hbda5;
mem_array[13783] = 16'ha28f;
mem_array[13782] = 16'h3da3;
mem_array[13785] = 16'hce98;
mem_array[13784] = 16'hbf95;
mem_array[13787] = 16'h6d56;
mem_array[13786] = 16'hbbeb;
mem_array[13789] = 16'h3eda;
mem_array[13788] = 16'hbeb8;
mem_array[13791] = 16'hcd88;
mem_array[13790] = 16'hbdc2;
mem_array[13793] = 16'hc26d;
mem_array[13792] = 16'hbe54;
mem_array[13795] = 16'hf42f;
mem_array[13794] = 16'hbf46;
mem_array[13797] = 16'h17eb;
mem_array[13796] = 16'h3eb6;
mem_array[13799] = 16'h260c;
mem_array[13798] = 16'h3f0a;
mem_array[13801] = 16'h5fad;
mem_array[13800] = 16'hbee9;
mem_array[13803] = 16'ha129;
mem_array[13802] = 16'hbe86;
mem_array[13805] = 16'hc427;
mem_array[13804] = 16'h3c6b;
mem_array[13807] = 16'h3fbc;
mem_array[13806] = 16'h3e21;
mem_array[13809] = 16'h4b0e;
mem_array[13808] = 16'hbe84;
mem_array[13811] = 16'h6c50;
mem_array[13810] = 16'hbeeb;
mem_array[13813] = 16'h1269;
mem_array[13812] = 16'h3e1b;
mem_array[13815] = 16'h2791;
mem_array[13814] = 16'hbda7;
mem_array[13817] = 16'h8463;
mem_array[13816] = 16'hbe4a;
mem_array[13819] = 16'h6e12;
mem_array[13818] = 16'h3cfe;
mem_array[13821] = 16'h71d4;
mem_array[13820] = 16'h3d45;
mem_array[13823] = 16'h3bb7;
mem_array[13822] = 16'h3d40;
mem_array[13825] = 16'hf089;
mem_array[13824] = 16'hbe25;
mem_array[13827] = 16'hce2f;
mem_array[13826] = 16'hbe6b;
mem_array[13829] = 16'h2422;
mem_array[13828] = 16'hbe77;
mem_array[13831] = 16'hfba1;
mem_array[13830] = 16'h3e39;
mem_array[13833] = 16'ha2f9;
mem_array[13832] = 16'hbf11;
mem_array[13835] = 16'h7644;
mem_array[13834] = 16'hbcbe;
mem_array[13837] = 16'h776e;
mem_array[13836] = 16'h3e43;
mem_array[13839] = 16'hedb2;
mem_array[13838] = 16'hbdc8;
mem_array[13841] = 16'hc982;
mem_array[13840] = 16'hbdf6;
mem_array[13843] = 16'hbfc2;
mem_array[13842] = 16'h3d95;
mem_array[13845] = 16'hf7bb;
mem_array[13844] = 16'hbfd5;
mem_array[13847] = 16'h308c;
mem_array[13846] = 16'hbee4;
mem_array[13849] = 16'hcce4;
mem_array[13848] = 16'hbe94;
mem_array[13851] = 16'hf769;
mem_array[13850] = 16'hbe04;
mem_array[13853] = 16'h2cb5;
mem_array[13852] = 16'hbdce;
mem_array[13855] = 16'hfede;
mem_array[13854] = 16'hbe06;
mem_array[13857] = 16'haa23;
mem_array[13856] = 16'h3f18;
mem_array[13859] = 16'h702f;
mem_array[13858] = 16'h3edc;
mem_array[13861] = 16'h27d0;
mem_array[13860] = 16'h3e45;
mem_array[13863] = 16'h89b4;
mem_array[13862] = 16'hbe6b;
mem_array[13865] = 16'h7130;
mem_array[13864] = 16'h3e81;
mem_array[13867] = 16'h0605;
mem_array[13866] = 16'hbcf0;
mem_array[13869] = 16'h4e64;
mem_array[13868] = 16'h3c8c;
mem_array[13871] = 16'hab30;
mem_array[13870] = 16'hbe6e;
mem_array[13873] = 16'h11f1;
mem_array[13872] = 16'hbdb5;
mem_array[13875] = 16'hf541;
mem_array[13874] = 16'hbf1a;
mem_array[13877] = 16'h0cf8;
mem_array[13876] = 16'h3e18;
mem_array[13879] = 16'hc4b6;
mem_array[13878] = 16'h3d8e;
mem_array[13881] = 16'h9e8c;
mem_array[13880] = 16'hbcf8;
mem_array[13883] = 16'h334f;
mem_array[13882] = 16'hbc53;
mem_array[13885] = 16'h7c2b;
mem_array[13884] = 16'h3db4;
mem_array[13887] = 16'hfe9c;
mem_array[13886] = 16'h3d92;
mem_array[13889] = 16'hdef0;
mem_array[13888] = 16'hbbcd;
mem_array[13891] = 16'h793a;
mem_array[13890] = 16'h3dae;
mem_array[13893] = 16'he9b5;
mem_array[13892] = 16'hbe10;
mem_array[13895] = 16'h8010;
mem_array[13894] = 16'h3d82;
mem_array[13897] = 16'h549f;
mem_array[13896] = 16'h3e7c;
mem_array[13899] = 16'h3985;
mem_array[13898] = 16'hbdb1;
mem_array[13901] = 16'h9a00;
mem_array[13900] = 16'h3e6e;
mem_array[13903] = 16'h325a;
mem_array[13902] = 16'hbd93;
mem_array[13905] = 16'hde34;
mem_array[13904] = 16'hbe8c;
mem_array[13907] = 16'hf56f;
mem_array[13906] = 16'hbe84;
mem_array[13909] = 16'h2024;
mem_array[13908] = 16'h3d7c;
mem_array[13911] = 16'h67f9;
mem_array[13910] = 16'h3e58;
mem_array[13913] = 16'h091d;
mem_array[13912] = 16'h3e4e;
mem_array[13915] = 16'h76d7;
mem_array[13914] = 16'h3e09;
mem_array[13917] = 16'h3ddd;
mem_array[13916] = 16'h3e14;
mem_array[13919] = 16'hfd72;
mem_array[13918] = 16'hbc63;
mem_array[13921] = 16'h7df7;
mem_array[13920] = 16'h3d91;
mem_array[13923] = 16'h21cb;
mem_array[13922] = 16'h3df7;
mem_array[13925] = 16'h830d;
mem_array[13924] = 16'h3dba;
mem_array[13927] = 16'hc9aa;
mem_array[13926] = 16'h3d63;
mem_array[13929] = 16'h5daf;
mem_array[13928] = 16'h3e87;
mem_array[13931] = 16'hc9db;
mem_array[13930] = 16'hbe90;
mem_array[13933] = 16'hc664;
mem_array[13932] = 16'hbe80;
mem_array[13935] = 16'h19ee;
mem_array[13934] = 16'hbe1c;
mem_array[13937] = 16'ha474;
mem_array[13936] = 16'hbe00;
mem_array[13939] = 16'ha346;
mem_array[13938] = 16'hbf62;
mem_array[13941] = 16'h2d2c;
mem_array[13940] = 16'h3c99;
mem_array[13943] = 16'hd7f8;
mem_array[13942] = 16'h3c7f;
mem_array[13945] = 16'h879d;
mem_array[13944] = 16'hbe49;
mem_array[13947] = 16'hbc67;
mem_array[13946] = 16'hbde7;
mem_array[13949] = 16'heec1;
mem_array[13948] = 16'h3e4c;
mem_array[13951] = 16'hb58c;
mem_array[13950] = 16'h3db8;
mem_array[13953] = 16'he0a8;
mem_array[13952] = 16'hbd8d;
mem_array[13955] = 16'h852c;
mem_array[13954] = 16'h3d8f;
mem_array[13957] = 16'hcd6e;
mem_array[13956] = 16'h3e83;
mem_array[13959] = 16'h8f52;
mem_array[13958] = 16'hbdd7;
mem_array[13961] = 16'h06a4;
mem_array[13960] = 16'h3d4d;
mem_array[13963] = 16'h101d;
mem_array[13962] = 16'h3e12;
mem_array[13965] = 16'h032b;
mem_array[13964] = 16'hbc93;
mem_array[13967] = 16'h7f6e;
mem_array[13966] = 16'hbea9;
mem_array[13969] = 16'h098c;
mem_array[13968] = 16'h3d67;
mem_array[13971] = 16'he655;
mem_array[13970] = 16'h3cfd;
mem_array[13973] = 16'hc0e1;
mem_array[13972] = 16'h3bf6;
mem_array[13975] = 16'h33bb;
mem_array[13974] = 16'hbe02;
mem_array[13977] = 16'h8bcb;
mem_array[13976] = 16'h3d5c;
mem_array[13979] = 16'hb24a;
mem_array[13978] = 16'hbf14;
mem_array[13981] = 16'h7814;
mem_array[13980] = 16'h3d05;
mem_array[13983] = 16'h3f70;
mem_array[13982] = 16'hbda7;
mem_array[13985] = 16'hdf48;
mem_array[13984] = 16'hbda9;
mem_array[13987] = 16'h1907;
mem_array[13986] = 16'hbe1b;
mem_array[13989] = 16'hedbf;
mem_array[13988] = 16'h3d81;
mem_array[13991] = 16'ha75f;
mem_array[13990] = 16'hbe0f;
mem_array[13993] = 16'h335f;
mem_array[13992] = 16'h3d5b;
mem_array[13995] = 16'hfad3;
mem_array[13994] = 16'hbf46;
mem_array[13997] = 16'h695d;
mem_array[13996] = 16'hbe2c;
mem_array[13999] = 16'h8a67;
mem_array[13998] = 16'hbf08;
mem_array[14001] = 16'h9e9f;
mem_array[14000] = 16'hbd37;
mem_array[14003] = 16'h0a0d;
mem_array[14002] = 16'hbd9f;
mem_array[14005] = 16'haa5b;
mem_array[14004] = 16'hbd97;
mem_array[14007] = 16'had49;
mem_array[14006] = 16'h3e28;
mem_array[14009] = 16'hb469;
mem_array[14008] = 16'h3e20;
mem_array[14011] = 16'h3e6f;
mem_array[14010] = 16'hbd07;
mem_array[14013] = 16'h3192;
mem_array[14012] = 16'h3eb3;
mem_array[14015] = 16'h6c22;
mem_array[14014] = 16'h3df3;
mem_array[14017] = 16'hc27f;
mem_array[14016] = 16'h3cba;
mem_array[14019] = 16'h21c9;
mem_array[14018] = 16'h3d26;
mem_array[14021] = 16'hfac0;
mem_array[14020] = 16'h3e07;
mem_array[14023] = 16'h636e;
mem_array[14022] = 16'h3dfb;
mem_array[14025] = 16'h82bf;
mem_array[14024] = 16'hbe03;
mem_array[14027] = 16'h3b28;
mem_array[14026] = 16'hbdf2;
mem_array[14029] = 16'h0eed;
mem_array[14028] = 16'h3e61;
mem_array[14031] = 16'h5f30;
mem_array[14030] = 16'h3e4c;
mem_array[14033] = 16'h3291;
mem_array[14032] = 16'hbe59;
mem_array[14035] = 16'h333d;
mem_array[14034] = 16'hbee2;
mem_array[14037] = 16'h1ce7;
mem_array[14036] = 16'h3c35;
mem_array[14039] = 16'hfb60;
mem_array[14038] = 16'hbef2;
mem_array[14041] = 16'h6c21;
mem_array[14040] = 16'hbe40;
mem_array[14043] = 16'h3a26;
mem_array[14042] = 16'h3e23;
mem_array[14045] = 16'ha03d;
mem_array[14044] = 16'h3db0;
mem_array[14047] = 16'h3127;
mem_array[14046] = 16'hbeac;
mem_array[14049] = 16'h9324;
mem_array[14048] = 16'hbe02;
mem_array[14051] = 16'hb0b9;
mem_array[14050] = 16'h3d98;
mem_array[14053] = 16'h5aa6;
mem_array[14052] = 16'h3eb7;
mem_array[14055] = 16'h620d;
mem_array[14054] = 16'hbf58;
mem_array[14057] = 16'h4f54;
mem_array[14056] = 16'h3df6;
mem_array[14059] = 16'hb596;
mem_array[14058] = 16'hbe3a;
mem_array[14061] = 16'h85b1;
mem_array[14060] = 16'hbe22;
mem_array[14063] = 16'he9e0;
mem_array[14062] = 16'h3d88;
mem_array[14065] = 16'h998b;
mem_array[14064] = 16'hbd92;
mem_array[14067] = 16'h66f9;
mem_array[14066] = 16'h3eec;
mem_array[14069] = 16'ha613;
mem_array[14068] = 16'hbd4c;
mem_array[14071] = 16'h2c53;
mem_array[14070] = 16'hbd54;
mem_array[14073] = 16'h33c3;
mem_array[14072] = 16'h3e5b;
mem_array[14075] = 16'h641d;
mem_array[14074] = 16'h3e05;
mem_array[14077] = 16'h16a5;
mem_array[14076] = 16'h3de8;
mem_array[14079] = 16'h0188;
mem_array[14078] = 16'hbe2a;
mem_array[14081] = 16'hc76b;
mem_array[14080] = 16'hbe5c;
mem_array[14083] = 16'h7860;
mem_array[14082] = 16'hbe4d;
mem_array[14085] = 16'h04b6;
mem_array[14084] = 16'hbf38;
mem_array[14087] = 16'hfc06;
mem_array[14086] = 16'hbdd3;
mem_array[14089] = 16'h5bfc;
mem_array[14088] = 16'h3e83;
mem_array[14091] = 16'hf5d4;
mem_array[14090] = 16'h3edd;
mem_array[14093] = 16'he3bb;
mem_array[14092] = 16'hbe22;
mem_array[14095] = 16'hfd3d;
mem_array[14094] = 16'hbed1;
mem_array[14097] = 16'h3ce7;
mem_array[14096] = 16'h3e38;
mem_array[14099] = 16'hc7ff;
mem_array[14098] = 16'hbecb;
mem_array[14101] = 16'h1f69;
mem_array[14100] = 16'hbf18;
mem_array[14103] = 16'hf010;
mem_array[14102] = 16'hbd1b;
mem_array[14105] = 16'h1975;
mem_array[14104] = 16'h3da7;
mem_array[14107] = 16'h7036;
mem_array[14106] = 16'hbdb5;
mem_array[14109] = 16'he6c3;
mem_array[14108] = 16'h3d35;
mem_array[14111] = 16'hf2df;
mem_array[14110] = 16'h3ebe;
mem_array[14113] = 16'h6bbc;
mem_array[14112] = 16'hbeb5;
mem_array[14115] = 16'h724b;
mem_array[14114] = 16'hbf8f;
mem_array[14117] = 16'h118b;
mem_array[14116] = 16'h3ddd;
mem_array[14119] = 16'h298c;
mem_array[14118] = 16'hbeab;
mem_array[14121] = 16'hd70c;
mem_array[14120] = 16'hbd02;
mem_array[14123] = 16'h468c;
mem_array[14122] = 16'hbcd8;
mem_array[14125] = 16'h2e57;
mem_array[14124] = 16'hbe94;
mem_array[14127] = 16'h8b5e;
mem_array[14126] = 16'hbe00;
mem_array[14129] = 16'hbe67;
mem_array[14128] = 16'hbd27;
mem_array[14131] = 16'h8905;
mem_array[14130] = 16'h3d83;
mem_array[14133] = 16'hbe27;
mem_array[14132] = 16'h3ed9;
mem_array[14135] = 16'hfa22;
mem_array[14134] = 16'h3c11;
mem_array[14137] = 16'h60b9;
mem_array[14136] = 16'h3e81;
mem_array[14139] = 16'hf89a;
mem_array[14138] = 16'hbdfd;
mem_array[14141] = 16'hde74;
mem_array[14140] = 16'hbe43;
mem_array[14143] = 16'h3942;
mem_array[14142] = 16'hbdd1;
mem_array[14145] = 16'h6c05;
mem_array[14144] = 16'hbee8;
mem_array[14147] = 16'h9903;
mem_array[14146] = 16'h3d9b;
mem_array[14149] = 16'h662d;
mem_array[14148] = 16'h3ee2;
mem_array[14151] = 16'h6cfe;
mem_array[14150] = 16'hbbc0;
mem_array[14153] = 16'h085e;
mem_array[14152] = 16'hbdc1;
mem_array[14155] = 16'h278f;
mem_array[14154] = 16'hbe5c;
mem_array[14157] = 16'hce83;
mem_array[14156] = 16'h3db2;
mem_array[14159] = 16'ha25a;
mem_array[14158] = 16'hbe95;
mem_array[14161] = 16'h657a;
mem_array[14160] = 16'hbf60;
mem_array[14163] = 16'h44c8;
mem_array[14162] = 16'h3da4;
mem_array[14165] = 16'h4914;
mem_array[14164] = 16'h3d39;
mem_array[14167] = 16'h4fb3;
mem_array[14166] = 16'hbd66;
mem_array[14169] = 16'h77b2;
mem_array[14168] = 16'h3c40;
mem_array[14171] = 16'h5c56;
mem_array[14170] = 16'h3e7e;
mem_array[14173] = 16'ha914;
mem_array[14172] = 16'hbddc;
mem_array[14175] = 16'h1b89;
mem_array[14174] = 16'hbec9;
mem_array[14177] = 16'h2691;
mem_array[14176] = 16'hbdd3;
mem_array[14179] = 16'h8110;
mem_array[14178] = 16'hbe9c;
mem_array[14181] = 16'hbdf6;
mem_array[14180] = 16'h3bc3;
mem_array[14183] = 16'h3924;
mem_array[14182] = 16'hbd2f;
mem_array[14185] = 16'h64b7;
mem_array[14184] = 16'hbe5d;
mem_array[14187] = 16'h4759;
mem_array[14186] = 16'hbe6c;
mem_array[14189] = 16'hcc0d;
mem_array[14188] = 16'hbe66;
mem_array[14191] = 16'h20be;
mem_array[14190] = 16'hbc67;
mem_array[14193] = 16'haaa9;
mem_array[14192] = 16'hbd6b;
mem_array[14195] = 16'h2306;
mem_array[14194] = 16'h3e72;
mem_array[14197] = 16'h5c24;
mem_array[14196] = 16'h3e47;
mem_array[14199] = 16'h0117;
mem_array[14198] = 16'h3e3d;
mem_array[14201] = 16'he18f;
mem_array[14200] = 16'hbdcc;
mem_array[14203] = 16'hd421;
mem_array[14202] = 16'h3dbf;
mem_array[14205] = 16'h3bd1;
mem_array[14204] = 16'hbe20;
mem_array[14207] = 16'he4b1;
mem_array[14206] = 16'hbda6;
mem_array[14209] = 16'h1fae;
mem_array[14208] = 16'h3dd8;
mem_array[14211] = 16'hfed7;
mem_array[14210] = 16'h3d89;
mem_array[14213] = 16'h9b41;
mem_array[14212] = 16'hb9fe;
mem_array[14215] = 16'h8c76;
mem_array[14214] = 16'h3b23;
mem_array[14217] = 16'h86e2;
mem_array[14216] = 16'h3d9d;
mem_array[14219] = 16'h1238;
mem_array[14218] = 16'hbe50;
mem_array[14221] = 16'h8f8d;
mem_array[14220] = 16'hbf54;
mem_array[14223] = 16'heeea;
mem_array[14222] = 16'hbe5a;
mem_array[14225] = 16'haf8f;
mem_array[14224] = 16'hbdf4;
mem_array[14227] = 16'h5908;
mem_array[14226] = 16'hbe13;
mem_array[14229] = 16'hb151;
mem_array[14228] = 16'h3e70;
mem_array[14231] = 16'h7bc3;
mem_array[14230] = 16'h3d26;
mem_array[14233] = 16'hca57;
mem_array[14232] = 16'h3dd2;
mem_array[14235] = 16'h0d1b;
mem_array[14234] = 16'hbf2a;
mem_array[14237] = 16'h5a62;
mem_array[14236] = 16'h3e26;
mem_array[14239] = 16'hc0fa;
mem_array[14238] = 16'h3e95;
mem_array[14241] = 16'h4beb;
mem_array[14240] = 16'h3c25;
mem_array[14243] = 16'h2211;
mem_array[14242] = 16'h3d96;
mem_array[14245] = 16'hc81e;
mem_array[14244] = 16'hbea1;
mem_array[14247] = 16'h0b1b;
mem_array[14246] = 16'hbc63;
mem_array[14249] = 16'h7d89;
mem_array[14248] = 16'hbe88;
mem_array[14251] = 16'hdc75;
mem_array[14250] = 16'hbca2;
mem_array[14253] = 16'habde;
mem_array[14252] = 16'hbd87;
mem_array[14255] = 16'h2df4;
mem_array[14254] = 16'hbea5;
mem_array[14257] = 16'hfc37;
mem_array[14256] = 16'hbe0d;
mem_array[14259] = 16'h27dd;
mem_array[14258] = 16'h3ea1;
mem_array[14261] = 16'h5d78;
mem_array[14260] = 16'hbe6c;
mem_array[14263] = 16'h5dca;
mem_array[14262] = 16'h3cb9;
mem_array[14265] = 16'hd55e;
mem_array[14264] = 16'hbe67;
mem_array[14267] = 16'h9665;
mem_array[14266] = 16'hbd34;
mem_array[14269] = 16'hc46e;
mem_array[14268] = 16'h3ddf;
mem_array[14271] = 16'h2708;
mem_array[14270] = 16'hbe19;
mem_array[14273] = 16'hde7e;
mem_array[14272] = 16'h3e81;
mem_array[14275] = 16'h4bef;
mem_array[14274] = 16'hbe21;
mem_array[14277] = 16'h7455;
mem_array[14276] = 16'h3eeb;
mem_array[14279] = 16'h254a;
mem_array[14278] = 16'hbc37;
mem_array[14281] = 16'hce55;
mem_array[14280] = 16'hbe7b;
mem_array[14283] = 16'h8f4f;
mem_array[14282] = 16'hbed8;
mem_array[14285] = 16'h3267;
mem_array[14284] = 16'h3e78;
mem_array[14287] = 16'h2822;
mem_array[14286] = 16'h3ea7;
mem_array[14289] = 16'hd785;
mem_array[14288] = 16'h3c99;
mem_array[14291] = 16'h7ca8;
mem_array[14290] = 16'hbe51;
mem_array[14293] = 16'h7cea;
mem_array[14292] = 16'hbe10;
mem_array[14295] = 16'hc6e9;
mem_array[14294] = 16'hbe82;
mem_array[14297] = 16'h5bf0;
mem_array[14296] = 16'h3e24;
mem_array[14299] = 16'h8799;
mem_array[14298] = 16'h3f01;
mem_array[14301] = 16'h69ec;
mem_array[14300] = 16'hbd3e;
mem_array[14303] = 16'h6d52;
mem_array[14302] = 16'hbca5;
mem_array[14305] = 16'h7811;
mem_array[14304] = 16'hbe6d;
mem_array[14307] = 16'ha84c;
mem_array[14306] = 16'h3e25;
mem_array[14309] = 16'hc471;
mem_array[14308] = 16'hbe92;
mem_array[14311] = 16'h7763;
mem_array[14310] = 16'hbe69;
mem_array[14313] = 16'hf8ae;
mem_array[14312] = 16'hbe13;
mem_array[14315] = 16'h07eb;
mem_array[14314] = 16'hbfb3;
mem_array[14317] = 16'heb55;
mem_array[14316] = 16'hbd51;
mem_array[14319] = 16'h1189;
mem_array[14318] = 16'hbe53;
mem_array[14321] = 16'h1362;
mem_array[14320] = 16'h3b8a;
mem_array[14323] = 16'h3a6e;
mem_array[14322] = 16'h3cc1;
mem_array[14325] = 16'hd503;
mem_array[14324] = 16'hbe2b;
mem_array[14327] = 16'h0d23;
mem_array[14326] = 16'hbebe;
mem_array[14329] = 16'hdfe3;
mem_array[14328] = 16'h3e70;
mem_array[14331] = 16'h9d67;
mem_array[14330] = 16'hbdbb;
mem_array[14333] = 16'h75ac;
mem_array[14332] = 16'h3dfb;
mem_array[14335] = 16'h07c1;
mem_array[14334] = 16'hbead;
mem_array[14337] = 16'h669a;
mem_array[14336] = 16'hbe1e;
mem_array[14339] = 16'hed82;
mem_array[14338] = 16'hbef6;
mem_array[14341] = 16'h3205;
mem_array[14340] = 16'h3d9a;
mem_array[14343] = 16'hca26;
mem_array[14342] = 16'hbe2c;
mem_array[14345] = 16'h951b;
mem_array[14344] = 16'h3e1e;
mem_array[14347] = 16'h55f5;
mem_array[14346] = 16'h3eb6;
mem_array[14349] = 16'h19df;
mem_array[14348] = 16'hbeb1;
mem_array[14351] = 16'h6541;
mem_array[14350] = 16'hbf06;
mem_array[14353] = 16'h83e0;
mem_array[14352] = 16'h3e17;
mem_array[14355] = 16'hf3cc;
mem_array[14354] = 16'hbcaf;
mem_array[14357] = 16'h3029;
mem_array[14356] = 16'h3d89;
mem_array[14359] = 16'hb836;
mem_array[14358] = 16'h3e47;
mem_array[14361] = 16'haede;
mem_array[14360] = 16'hbd33;
mem_array[14363] = 16'hfcd1;
mem_array[14362] = 16'hbcb9;
mem_array[14365] = 16'h6d25;
mem_array[14364] = 16'hbe95;
mem_array[14367] = 16'h8939;
mem_array[14366] = 16'hbd2a;
mem_array[14369] = 16'h8559;
mem_array[14368] = 16'hbe87;
mem_array[14371] = 16'hb7b4;
mem_array[14370] = 16'hbd4f;
mem_array[14373] = 16'h4314;
mem_array[14372] = 16'hbeee;
mem_array[14375] = 16'h7eb9;
mem_array[14374] = 16'hbf1d;
mem_array[14377] = 16'he522;
mem_array[14376] = 16'h3e43;
mem_array[14379] = 16'hf7f7;
mem_array[14378] = 16'hbed3;
mem_array[14381] = 16'hd090;
mem_array[14380] = 16'h3ded;
mem_array[14383] = 16'h59ca;
mem_array[14382] = 16'h3e5b;
mem_array[14385] = 16'h053e;
mem_array[14384] = 16'hbe91;
mem_array[14387] = 16'h4e03;
mem_array[14386] = 16'hbe56;
mem_array[14389] = 16'hd2f2;
mem_array[14388] = 16'h3e6e;
mem_array[14391] = 16'h6d2b;
mem_array[14390] = 16'h3e39;
mem_array[14393] = 16'h40c9;
mem_array[14392] = 16'hbca7;
mem_array[14395] = 16'h02ad;
mem_array[14394] = 16'hbe26;
mem_array[14397] = 16'he9bc;
mem_array[14396] = 16'hbe93;
mem_array[14399] = 16'h89cf;
mem_array[14398] = 16'hbf03;
mem_array[14401] = 16'hc920;
mem_array[14400] = 16'h3e8f;
mem_array[14403] = 16'hcc0f;
mem_array[14402] = 16'h3dbf;
mem_array[14405] = 16'hde12;
mem_array[14404] = 16'hbd6c;
mem_array[14407] = 16'h6f84;
mem_array[14406] = 16'h3f1d;
mem_array[14409] = 16'h16ab;
mem_array[14408] = 16'hbe9a;
mem_array[14411] = 16'h59cc;
mem_array[14410] = 16'hbe69;
mem_array[14413] = 16'h93c6;
mem_array[14412] = 16'h3d9c;
mem_array[14415] = 16'h1ba1;
mem_array[14414] = 16'hbd7a;
mem_array[14417] = 16'h2648;
mem_array[14416] = 16'hbe92;
mem_array[14419] = 16'h55f9;
mem_array[14418] = 16'h3d5a;
mem_array[14421] = 16'h7771;
mem_array[14420] = 16'hbde1;
mem_array[14423] = 16'hb20b;
mem_array[14422] = 16'h3ccd;
mem_array[14425] = 16'h654d;
mem_array[14424] = 16'hbe1b;
mem_array[14427] = 16'h2dc1;
mem_array[14426] = 16'h3d6e;
mem_array[14429] = 16'h958e;
mem_array[14428] = 16'hbe97;
mem_array[14431] = 16'hcb10;
mem_array[14430] = 16'hbe42;
mem_array[14433] = 16'hd249;
mem_array[14432] = 16'hbd7c;
mem_array[14435] = 16'hcef2;
mem_array[14434] = 16'h3e34;
mem_array[14437] = 16'hac69;
mem_array[14436] = 16'h3cd7;
mem_array[14439] = 16'h7cd5;
mem_array[14438] = 16'hbf07;
mem_array[14441] = 16'h29c7;
mem_array[14440] = 16'hbeb7;
mem_array[14443] = 16'h2028;
mem_array[14442] = 16'h3e81;
mem_array[14445] = 16'h002e;
mem_array[14444] = 16'hbe0d;
mem_array[14447] = 16'hfdfa;
mem_array[14446] = 16'hbcd2;
mem_array[14449] = 16'hf1b7;
mem_array[14448] = 16'hbdfe;
mem_array[14451] = 16'h211a;
mem_array[14450] = 16'h3da5;
mem_array[14453] = 16'hc3d4;
mem_array[14452] = 16'hbdaf;
mem_array[14455] = 16'h1cbc;
mem_array[14454] = 16'hbd81;
mem_array[14457] = 16'hdb83;
mem_array[14456] = 16'hbe38;
mem_array[14459] = 16'h0d3f;
mem_array[14458] = 16'hbf03;
mem_array[14461] = 16'hb84c;
mem_array[14460] = 16'h3edc;
mem_array[14463] = 16'h69f3;
mem_array[14462] = 16'hbdcb;
mem_array[14465] = 16'hf442;
mem_array[14464] = 16'hbe84;
mem_array[14467] = 16'h8d02;
mem_array[14466] = 16'h3ef0;
mem_array[14469] = 16'h34cb;
mem_array[14468] = 16'hbe78;
mem_array[14471] = 16'h880b;
mem_array[14470] = 16'hbe3d;
mem_array[14473] = 16'hd6dc;
mem_array[14472] = 16'h3cf7;
mem_array[14475] = 16'he09c;
mem_array[14474] = 16'hbd7b;
mem_array[14477] = 16'h2ddf;
mem_array[14476] = 16'hbeda;
mem_array[14479] = 16'h76b5;
mem_array[14478] = 16'hbd68;
mem_array[14481] = 16'h79a1;
mem_array[14480] = 16'hbdc1;
mem_array[14483] = 16'hb753;
mem_array[14482] = 16'hbd9a;
mem_array[14485] = 16'haee0;
mem_array[14484] = 16'hbe33;
mem_array[14487] = 16'hff2e;
mem_array[14486] = 16'hbd08;
mem_array[14489] = 16'h784f;
mem_array[14488] = 16'hbe73;
mem_array[14491] = 16'hbfbd;
mem_array[14490] = 16'hbc93;
mem_array[14493] = 16'hcfd9;
mem_array[14492] = 16'h3e9e;
mem_array[14495] = 16'hf3dd;
mem_array[14494] = 16'h3eac;
mem_array[14497] = 16'hadae;
mem_array[14496] = 16'h3e25;
mem_array[14499] = 16'h97ec;
mem_array[14498] = 16'hbe6b;
mem_array[14501] = 16'hbc82;
mem_array[14500] = 16'hbe5d;
mem_array[14503] = 16'h2a24;
mem_array[14502] = 16'h3e6b;
mem_array[14505] = 16'h9c9b;
mem_array[14504] = 16'hbd77;
mem_array[14507] = 16'h30d0;
mem_array[14506] = 16'h3d38;
mem_array[14509] = 16'h289e;
mem_array[14508] = 16'h3d89;
mem_array[14511] = 16'h2349;
mem_array[14510] = 16'h3e0a;
mem_array[14513] = 16'h1a81;
mem_array[14512] = 16'hbe85;
mem_array[14515] = 16'hc46b;
mem_array[14514] = 16'hbd72;
mem_array[14517] = 16'h34cc;
mem_array[14516] = 16'hbd5e;
mem_array[14519] = 16'h588e;
mem_array[14518] = 16'hbe76;
mem_array[14521] = 16'h9030;
mem_array[14520] = 16'hbd90;
mem_array[14523] = 16'hdcd4;
mem_array[14522] = 16'h3aa9;
mem_array[14525] = 16'hab31;
mem_array[14524] = 16'h3cc6;
mem_array[14527] = 16'hd839;
mem_array[14526] = 16'h3eb2;
mem_array[14529] = 16'h0794;
mem_array[14528] = 16'h3e78;
mem_array[14531] = 16'h7f1c;
mem_array[14530] = 16'h3ee9;
mem_array[14533] = 16'ha5a2;
mem_array[14532] = 16'hbd30;
mem_array[14535] = 16'hc8d6;
mem_array[14534] = 16'h3e24;
mem_array[14537] = 16'h751b;
mem_array[14536] = 16'hbe64;
mem_array[14539] = 16'hc0d0;
mem_array[14538] = 16'hbe14;
mem_array[14541] = 16'h6c45;
mem_array[14540] = 16'hbd49;
mem_array[14543] = 16'h5b0a;
mem_array[14542] = 16'h3d62;
mem_array[14545] = 16'hcc83;
mem_array[14544] = 16'hbe5f;
mem_array[14547] = 16'h3e0e;
mem_array[14546] = 16'hbcde;
mem_array[14549] = 16'he3c6;
mem_array[14548] = 16'h3e92;
mem_array[14551] = 16'hea0e;
mem_array[14550] = 16'hbe09;
mem_array[14553] = 16'h4f8b;
mem_array[14552] = 16'hbc3e;
mem_array[14555] = 16'he69f;
mem_array[14554] = 16'h3d98;
mem_array[14557] = 16'h2f65;
mem_array[14556] = 16'h3e62;
mem_array[14559] = 16'hddb4;
mem_array[14558] = 16'hbcb1;
mem_array[14561] = 16'h01e7;
mem_array[14560] = 16'hbe20;
mem_array[14563] = 16'h903c;
mem_array[14562] = 16'hbd84;
mem_array[14565] = 16'hb988;
mem_array[14564] = 16'hbf2b;
mem_array[14567] = 16'ha482;
mem_array[14566] = 16'hbe22;
mem_array[14569] = 16'h7e3a;
mem_array[14568] = 16'h3dd7;
mem_array[14571] = 16'h7f2b;
mem_array[14570] = 16'h3ed1;
mem_array[14573] = 16'h05ba;
mem_array[14572] = 16'h3d92;
mem_array[14575] = 16'h0c69;
mem_array[14574] = 16'hbdc7;
mem_array[14577] = 16'h9c4d;
mem_array[14576] = 16'hbe68;
mem_array[14579] = 16'h0f4e;
mem_array[14578] = 16'hbef9;
mem_array[14581] = 16'h2484;
mem_array[14580] = 16'hbd3d;
mem_array[14583] = 16'h172d;
mem_array[14582] = 16'hbe84;
mem_array[14585] = 16'hd729;
mem_array[14584] = 16'hbd85;
mem_array[14587] = 16'hf2d7;
mem_array[14586] = 16'h3e01;
mem_array[14589] = 16'hf453;
mem_array[14588] = 16'h3e97;
mem_array[14591] = 16'h1d11;
mem_array[14590] = 16'h3e9e;
mem_array[14593] = 16'h8f62;
mem_array[14592] = 16'h3e27;
mem_array[14595] = 16'ha818;
mem_array[14594] = 16'hbced;
mem_array[14597] = 16'hf870;
mem_array[14596] = 16'h3e70;
mem_array[14599] = 16'h3f55;
mem_array[14598] = 16'hbe04;
mem_array[14601] = 16'heda5;
mem_array[14600] = 16'h3c35;
mem_array[14603] = 16'h2570;
mem_array[14602] = 16'hbbcc;
mem_array[14605] = 16'hf44c;
mem_array[14604] = 16'hbda1;
mem_array[14607] = 16'h3332;
mem_array[14606] = 16'h3d9d;
mem_array[14609] = 16'hb302;
mem_array[14608] = 16'h3e99;
mem_array[14611] = 16'h1ca7;
mem_array[14610] = 16'h3d7c;
mem_array[14613] = 16'h9eec;
mem_array[14612] = 16'h3d07;
mem_array[14615] = 16'hf8f1;
mem_array[14614] = 16'hbcb6;
mem_array[14617] = 16'hac1d;
mem_array[14616] = 16'hbd40;
mem_array[14619] = 16'h1b4d;
mem_array[14618] = 16'hbde9;
mem_array[14621] = 16'hef91;
mem_array[14620] = 16'hbeac;
mem_array[14623] = 16'h99fc;
mem_array[14622] = 16'hbcac;
mem_array[14625] = 16'h172a;
mem_array[14624] = 16'hbfe0;
mem_array[14627] = 16'h39d1;
mem_array[14626] = 16'h3c8f;
mem_array[14629] = 16'ha1b9;
mem_array[14628] = 16'h3e24;
mem_array[14631] = 16'h6323;
mem_array[14630] = 16'h3e4f;
mem_array[14633] = 16'h67ad;
mem_array[14632] = 16'h3e3f;
mem_array[14635] = 16'hb4d7;
mem_array[14634] = 16'h3d78;
mem_array[14637] = 16'hdcbc;
mem_array[14636] = 16'hbe40;
mem_array[14639] = 16'he799;
mem_array[14638] = 16'hbef9;
mem_array[14641] = 16'h3584;
mem_array[14640] = 16'h3ccf;
mem_array[14643] = 16'haca2;
mem_array[14642] = 16'hbf0d;
mem_array[14645] = 16'hc08c;
mem_array[14644] = 16'hbe7e;
mem_array[14647] = 16'hfdc4;
mem_array[14646] = 16'h3e07;
mem_array[14649] = 16'h8b18;
mem_array[14648] = 16'h3def;
mem_array[14651] = 16'h5b12;
mem_array[14650] = 16'h3f11;
mem_array[14653] = 16'h20d4;
mem_array[14652] = 16'h3d31;
mem_array[14655] = 16'h9cda;
mem_array[14654] = 16'h3da0;
mem_array[14657] = 16'ha29c;
mem_array[14656] = 16'h3d58;
mem_array[14659] = 16'hf834;
mem_array[14658] = 16'hbf87;
mem_array[14661] = 16'h05ba;
mem_array[14660] = 16'hbdb9;
mem_array[14663] = 16'hc429;
mem_array[14662] = 16'hbd82;
mem_array[14665] = 16'hf352;
mem_array[14664] = 16'hbe20;
mem_array[14667] = 16'h43f7;
mem_array[14666] = 16'hbe9f;
mem_array[14669] = 16'hdc3f;
mem_array[14668] = 16'h3e1b;
mem_array[14671] = 16'h5be3;
mem_array[14670] = 16'h3cb3;
mem_array[14673] = 16'h92c0;
mem_array[14672] = 16'hbde2;
mem_array[14675] = 16'h4295;
mem_array[14674] = 16'hbd92;
mem_array[14677] = 16'he33d;
mem_array[14676] = 16'hbe4a;
mem_array[14679] = 16'ha063;
mem_array[14678] = 16'h3dd6;
mem_array[14681] = 16'hbe05;
mem_array[14680] = 16'hbe81;
mem_array[14683] = 16'h2985;
mem_array[14682] = 16'h3c58;
mem_array[14685] = 16'h9e27;
mem_array[14684] = 16'hbfe8;
mem_array[14687] = 16'hc0b9;
mem_array[14686] = 16'hbcb2;
mem_array[14689] = 16'h6d3e;
mem_array[14688] = 16'hbdc4;
mem_array[14691] = 16'hf381;
mem_array[14690] = 16'hbe04;
mem_array[14693] = 16'hcadb;
mem_array[14692] = 16'h3e05;
mem_array[14695] = 16'hfc9a;
mem_array[14694] = 16'h3e27;
mem_array[14697] = 16'h3b2d;
mem_array[14696] = 16'hbdac;
mem_array[14699] = 16'h1a2b;
mem_array[14698] = 16'hbdde;
mem_array[14701] = 16'hde7d;
mem_array[14700] = 16'hbe4a;
mem_array[14703] = 16'he974;
mem_array[14702] = 16'h3e45;
mem_array[14705] = 16'h6953;
mem_array[14704] = 16'hbe95;
mem_array[14707] = 16'he3fd;
mem_array[14706] = 16'hbe18;
mem_array[14709] = 16'h45d8;
mem_array[14708] = 16'hbdf1;
mem_array[14711] = 16'h60af;
mem_array[14710] = 16'h3f17;
mem_array[14713] = 16'h676f;
mem_array[14712] = 16'h3e93;
mem_array[14715] = 16'h3cfb;
mem_array[14714] = 16'h3d33;
mem_array[14717] = 16'h1c94;
mem_array[14716] = 16'hbe40;
mem_array[14719] = 16'h77d3;
mem_array[14718] = 16'hbdf9;
mem_array[14721] = 16'h23e2;
mem_array[14720] = 16'hbd6d;
mem_array[14723] = 16'hfcea;
mem_array[14722] = 16'hbdcf;
mem_array[14725] = 16'h4d2f;
mem_array[14724] = 16'h3d97;
mem_array[14727] = 16'h394c;
mem_array[14726] = 16'hbdfa;
mem_array[14729] = 16'hd237;
mem_array[14728] = 16'hbcb2;
mem_array[14731] = 16'h2491;
mem_array[14730] = 16'h3d52;
mem_array[14733] = 16'h7711;
mem_array[14732] = 16'h3d8e;
mem_array[14735] = 16'h7dbd;
mem_array[14734] = 16'h3ddb;
mem_array[14737] = 16'h8095;
mem_array[14736] = 16'hbbf5;
mem_array[14739] = 16'h05d2;
mem_array[14738] = 16'h3ebb;
mem_array[14741] = 16'h308f;
mem_array[14740] = 16'hbd89;
mem_array[14743] = 16'h4056;
mem_array[14742] = 16'hbd86;
mem_array[14745] = 16'h6d69;
mem_array[14744] = 16'hbf3b;
mem_array[14747] = 16'h9e80;
mem_array[14746] = 16'hbd09;
mem_array[14749] = 16'hc56a;
mem_array[14748] = 16'h3d44;
mem_array[14751] = 16'hd398;
mem_array[14750] = 16'h3ea4;
mem_array[14753] = 16'h8566;
mem_array[14752] = 16'hbe1d;
mem_array[14755] = 16'h7785;
mem_array[14754] = 16'h3a6f;
mem_array[14757] = 16'h76d9;
mem_array[14756] = 16'hbe39;
mem_array[14759] = 16'ha0b7;
mem_array[14758] = 16'hbce9;
mem_array[14761] = 16'hba3b;
mem_array[14760] = 16'hbebf;
mem_array[14763] = 16'h7069;
mem_array[14762] = 16'hbdfa;
mem_array[14765] = 16'h0e1e;
mem_array[14764] = 16'hbdb5;
mem_array[14767] = 16'h0255;
mem_array[14766] = 16'h3d54;
mem_array[14769] = 16'h1d09;
mem_array[14768] = 16'hbd0a;
mem_array[14771] = 16'he845;
mem_array[14770] = 16'h3e9b;
mem_array[14773] = 16'h460b;
mem_array[14772] = 16'hbe85;
mem_array[14775] = 16'hb563;
mem_array[14774] = 16'h3e9c;
mem_array[14777] = 16'h129c;
mem_array[14776] = 16'hbcb7;
mem_array[14779] = 16'hb1ab;
mem_array[14778] = 16'hbdad;
mem_array[14781] = 16'h12cd;
mem_array[14780] = 16'hbc33;
mem_array[14783] = 16'hcd2b;
mem_array[14782] = 16'hbc72;
mem_array[14785] = 16'h9127;
mem_array[14784] = 16'hbe86;
mem_array[14787] = 16'hf3b1;
mem_array[14786] = 16'h3e6a;
mem_array[14789] = 16'h7f57;
mem_array[14788] = 16'h3cc5;
mem_array[14791] = 16'h5301;
mem_array[14790] = 16'h3e17;
mem_array[14793] = 16'hf33f;
mem_array[14792] = 16'hbec5;
mem_array[14795] = 16'h4d91;
mem_array[14794] = 16'h3ea6;
mem_array[14797] = 16'h025a;
mem_array[14796] = 16'hbe9b;
mem_array[14799] = 16'h28b9;
mem_array[14798] = 16'hbc9b;
mem_array[14801] = 16'hd29d;
mem_array[14800] = 16'h3e16;
mem_array[14803] = 16'hac66;
mem_array[14802] = 16'h3e32;
mem_array[14805] = 16'h4842;
mem_array[14804] = 16'hbe47;
mem_array[14807] = 16'h452a;
mem_array[14806] = 16'hbe1d;
mem_array[14809] = 16'hf7da;
mem_array[14808] = 16'h3dbd;
mem_array[14811] = 16'h4f6b;
mem_array[14810] = 16'hbe83;
mem_array[14813] = 16'hc751;
mem_array[14812] = 16'h3e9b;
mem_array[14815] = 16'h842b;
mem_array[14814] = 16'h3e30;
mem_array[14817] = 16'h5182;
mem_array[14816] = 16'hbeb9;
mem_array[14819] = 16'h8624;
mem_array[14818] = 16'h3e37;
mem_array[14821] = 16'hc926;
mem_array[14820] = 16'hbe73;
mem_array[14823] = 16'hf31b;
mem_array[14822] = 16'h3cba;
mem_array[14825] = 16'hd053;
mem_array[14824] = 16'h3eb8;
mem_array[14827] = 16'h9f11;
mem_array[14826] = 16'h3eab;
mem_array[14829] = 16'h7fca;
mem_array[14828] = 16'h3dad;
mem_array[14831] = 16'h9e14;
mem_array[14830] = 16'h3ec0;
mem_array[14833] = 16'he412;
mem_array[14832] = 16'hc02e;
mem_array[14835] = 16'h6db8;
mem_array[14834] = 16'hbba5;
mem_array[14837] = 16'h94a4;
mem_array[14836] = 16'hbf28;
mem_array[14839] = 16'hdf6a;
mem_array[14838] = 16'h3de9;
mem_array[14841] = 16'h5fce;
mem_array[14840] = 16'h3d30;
mem_array[14843] = 16'h177a;
mem_array[14842] = 16'h3cc4;
mem_array[14845] = 16'ha6d1;
mem_array[14844] = 16'hbeaf;
mem_array[14847] = 16'h9481;
mem_array[14846] = 16'hbeff;
mem_array[14849] = 16'h46cc;
mem_array[14848] = 16'h3e87;
mem_array[14851] = 16'h8483;
mem_array[14850] = 16'hbccd;
mem_array[14853] = 16'hbb24;
mem_array[14852] = 16'hbe88;
mem_array[14855] = 16'h1a0c;
mem_array[14854] = 16'h3e2d;
mem_array[14857] = 16'h15cf;
mem_array[14856] = 16'hbf4e;
mem_array[14859] = 16'h2cd6;
mem_array[14858] = 16'h3ead;
mem_array[14861] = 16'hde4f;
mem_array[14860] = 16'h3cd8;
mem_array[14863] = 16'h26ed;
mem_array[14862] = 16'h3e91;
mem_array[14865] = 16'h68e6;
mem_array[14864] = 16'hbf4d;
mem_array[14867] = 16'h4a64;
mem_array[14866] = 16'hbe0f;
mem_array[14869] = 16'h02f9;
mem_array[14868] = 16'hbf09;
mem_array[14871] = 16'h716e;
mem_array[14870] = 16'h3ddc;
mem_array[14873] = 16'h6a06;
mem_array[14872] = 16'h3f0a;
mem_array[14875] = 16'ha804;
mem_array[14874] = 16'h3e88;
mem_array[14877] = 16'h3bc5;
mem_array[14876] = 16'hbfa0;
mem_array[14879] = 16'h5007;
mem_array[14878] = 16'hbf46;
mem_array[14881] = 16'h6f95;
mem_array[14880] = 16'hbf9c;
mem_array[14883] = 16'h8f77;
mem_array[14882] = 16'hbd80;
mem_array[14885] = 16'hf6e8;
mem_array[14884] = 16'hbe95;
mem_array[14887] = 16'haeb6;
mem_array[14886] = 16'hbe93;
mem_array[14889] = 16'hb71d;
mem_array[14888] = 16'hbd9f;
mem_array[14891] = 16'hc366;
mem_array[14890] = 16'h3e91;
mem_array[14893] = 16'h1ba3;
mem_array[14892] = 16'hc03f;
mem_array[14895] = 16'h6e50;
mem_array[14894] = 16'h3ea3;
mem_array[14897] = 16'he5cb;
mem_array[14896] = 16'hbfcd;
mem_array[14899] = 16'h4b3f;
mem_array[14898] = 16'hbf63;
mem_array[14901] = 16'hc60b;
mem_array[14900] = 16'h3d99;
mem_array[14903] = 16'h42c7;
mem_array[14902] = 16'h3dae;
mem_array[14905] = 16'h275c;
mem_array[14904] = 16'hbfc1;
mem_array[14907] = 16'he1bf;
mem_array[14906] = 16'hbf79;
mem_array[14909] = 16'hb7ed;
mem_array[14908] = 16'hbfb2;
mem_array[14911] = 16'hf4d3;
mem_array[14910] = 16'hbe90;
mem_array[14913] = 16'h5fd3;
mem_array[14912] = 16'hbf48;
mem_array[14915] = 16'h13ab;
mem_array[14914] = 16'hbf07;
mem_array[14917] = 16'h3bf0;
mem_array[14916] = 16'hbfab;
mem_array[14919] = 16'hf3a2;
mem_array[14918] = 16'h3eef;
mem_array[14921] = 16'h42f9;
mem_array[14920] = 16'h3eb7;
mem_array[14923] = 16'hab1f;
mem_array[14922] = 16'hbc1e;
mem_array[14925] = 16'h5909;
mem_array[14924] = 16'hbf52;
mem_array[14927] = 16'h4c5e;
mem_array[14926] = 16'hbe6b;
mem_array[14929] = 16'hca15;
mem_array[14928] = 16'hbfa9;
mem_array[14931] = 16'h0e6b;
mem_array[14930] = 16'h3e6b;
mem_array[14933] = 16'h2fa8;
mem_array[14932] = 16'h3f28;
mem_array[14935] = 16'h6d75;
mem_array[14934] = 16'h3f3c;
mem_array[14937] = 16'hf312;
mem_array[14936] = 16'hbfa9;
mem_array[14939] = 16'hbe10;
mem_array[14938] = 16'hbf64;
mem_array[14941] = 16'h0aa3;
mem_array[14940] = 16'hbfd4;
mem_array[14943] = 16'h31ad;
mem_array[14942] = 16'hbec0;
mem_array[14945] = 16'hbb21;
mem_array[14944] = 16'hbf62;
mem_array[14947] = 16'hee8a;
mem_array[14946] = 16'hbfdc;
mem_array[14949] = 16'h555b;
mem_array[14948] = 16'h3f2d;
mem_array[14951] = 16'h081b;
mem_array[14950] = 16'h3ea5;
mem_array[14953] = 16'h95c0;
mem_array[14952] = 16'hbfd6;
mem_array[14955] = 16'h2bf8;
mem_array[14954] = 16'h3eaf;
mem_array[14957] = 16'h39c8;
mem_array[14956] = 16'hbf6b;
mem_array[14959] = 16'hf882;
mem_array[14958] = 16'hbf32;
mem_array[14961] = 16'h10a6;
mem_array[14960] = 16'hbddd;
mem_array[14963] = 16'hbccb;
mem_array[14962] = 16'hbd50;
mem_array[14965] = 16'h0165;
mem_array[14964] = 16'hbfcd;
mem_array[14967] = 16'h980b;
mem_array[14966] = 16'h3e9c;
mem_array[14969] = 16'h8d43;
mem_array[14968] = 16'hbf48;
mem_array[14971] = 16'h10a2;
mem_array[14970] = 16'hbea0;
mem_array[14973] = 16'h1575;
mem_array[14972] = 16'hbf9b;
mem_array[14975] = 16'h7dd9;
mem_array[14974] = 16'h3e99;
mem_array[14977] = 16'h8d6f;
mem_array[14976] = 16'hbfb3;
mem_array[14979] = 16'h1fed;
mem_array[14978] = 16'h3e77;
mem_array[14981] = 16'hbdc5;
mem_array[14980] = 16'h3f03;
mem_array[14983] = 16'hfd48;
mem_array[14982] = 16'h3d6a;
mem_array[14985] = 16'h31db;
mem_array[14984] = 16'hbef5;
mem_array[14987] = 16'h7090;
mem_array[14986] = 16'hbe6c;
mem_array[14989] = 16'h2784;
mem_array[14988] = 16'hbf8f;
mem_array[14991] = 16'habb6;
mem_array[14990] = 16'hbf51;
mem_array[14993] = 16'h353f;
mem_array[14992] = 16'h3eae;
mem_array[14995] = 16'h953f;
mem_array[14994] = 16'h3ec7;
mem_array[14997] = 16'h29d4;
mem_array[14996] = 16'hbe8b;
mem_array[14999] = 16'h9e0f;
mem_array[14998] = 16'hbf9f;
mem_array[15001] = 16'h886c;
mem_array[15000] = 16'h3dc3;
mem_array[15003] = 16'h7391;
mem_array[15002] = 16'hbf54;
mem_array[15005] = 16'h7b14;
mem_array[15004] = 16'hbe98;
mem_array[15007] = 16'h682f;
mem_array[15006] = 16'hbfe3;
mem_array[15009] = 16'hefb7;
mem_array[15008] = 16'h3eeb;
mem_array[15011] = 16'hb962;
mem_array[15010] = 16'h3ead;
mem_array[15013] = 16'h3c4c;
mem_array[15012] = 16'hbf0e;
mem_array[15015] = 16'h82f9;
mem_array[15014] = 16'h3dda;
mem_array[15017] = 16'h8d9d;
mem_array[15016] = 16'hbdd3;
mem_array[15019] = 16'habd7;
mem_array[15018] = 16'h3ea0;
mem_array[15021] = 16'he31c;
mem_array[15020] = 16'h3c86;
mem_array[15023] = 16'ha319;
mem_array[15022] = 16'hbb9e;
mem_array[15025] = 16'h1b51;
mem_array[15024] = 16'hbf1d;
mem_array[15027] = 16'head5;
mem_array[15026] = 16'hbd21;
mem_array[15029] = 16'hfac9;
mem_array[15028] = 16'hbf42;
mem_array[15031] = 16'hf9cb;
mem_array[15030] = 16'h3e11;
mem_array[15033] = 16'hdc4f;
mem_array[15032] = 16'h3d54;
mem_array[15035] = 16'h30be;
mem_array[15034] = 16'hbfc9;
mem_array[15037] = 16'h8996;
mem_array[15036] = 16'hbee1;
mem_array[15039] = 16'hcde0;
mem_array[15038] = 16'hbe64;
mem_array[15041] = 16'hc988;
mem_array[15040] = 16'hbe8e;
mem_array[15043] = 16'ha63a;
mem_array[15042] = 16'hbf22;
mem_array[15045] = 16'h88ea;
mem_array[15044] = 16'hbe42;
mem_array[15047] = 16'haf69;
mem_array[15046] = 16'hbf26;
mem_array[15049] = 16'h8b14;
mem_array[15048] = 16'hbf8a;
mem_array[15051] = 16'h4e0d;
mem_array[15050] = 16'hbf09;
mem_array[15053] = 16'h6d0f;
mem_array[15052] = 16'h3e9d;
mem_array[15055] = 16'hf04c;
mem_array[15054] = 16'h3e6e;
mem_array[15057] = 16'h02cf;
mem_array[15056] = 16'hbc31;
mem_array[15059] = 16'h0f8a;
mem_array[15058] = 16'hbf8f;
mem_array[15061] = 16'h9f77;
mem_array[15060] = 16'h3e25;
mem_array[15063] = 16'hd27a;
mem_array[15062] = 16'hbf06;
mem_array[15065] = 16'h7c8e;
mem_array[15064] = 16'hbe63;
mem_array[15067] = 16'hb365;
mem_array[15066] = 16'hbe99;
mem_array[15069] = 16'h3c4a;
mem_array[15068] = 16'hbd99;
mem_array[15071] = 16'h401b;
mem_array[15070] = 16'h3f22;
mem_array[15073] = 16'hb71f;
mem_array[15072] = 16'h3e77;
mem_array[15075] = 16'h34ec;
mem_array[15074] = 16'hbf34;
mem_array[15077] = 16'h674f;
mem_array[15076] = 16'hbd7b;
mem_array[15079] = 16'h88bf;
mem_array[15078] = 16'h3db7;
mem_array[15081] = 16'h3564;
mem_array[15080] = 16'h3a92;
mem_array[15083] = 16'hb56c;
mem_array[15082] = 16'hbb64;
mem_array[15085] = 16'h82f5;
mem_array[15084] = 16'hbe24;
mem_array[15087] = 16'h3ca0;
mem_array[15086] = 16'hbc64;
mem_array[15089] = 16'h1a2f;
mem_array[15088] = 16'hbdb9;
mem_array[15091] = 16'h42aa;
mem_array[15090] = 16'h3f56;
mem_array[15093] = 16'hb8b7;
mem_array[15092] = 16'h3d44;
mem_array[15095] = 16'h1b96;
mem_array[15094] = 16'hbf6f;
mem_array[15097] = 16'hd0d4;
mem_array[15096] = 16'hbf20;
mem_array[15099] = 16'hd90d;
mem_array[15098] = 16'hbf67;
mem_array[15101] = 16'h43de;
mem_array[15100] = 16'hbef1;
mem_array[15103] = 16'h94bf;
mem_array[15102] = 16'hbf63;
mem_array[15105] = 16'h978a;
mem_array[15104] = 16'hbd92;
mem_array[15107] = 16'hcd8e;
mem_array[15106] = 16'hbeb7;
mem_array[15109] = 16'ha9fd;
mem_array[15108] = 16'hbd96;
mem_array[15111] = 16'hd62f;
mem_array[15110] = 16'hbebe;
mem_array[15113] = 16'h0eef;
mem_array[15112] = 16'h3cf2;
mem_array[15115] = 16'h540d;
mem_array[15114] = 16'h3e86;
mem_array[15117] = 16'hbed7;
mem_array[15116] = 16'h3dcd;
mem_array[15119] = 16'hba61;
mem_array[15118] = 16'h3d9d;
mem_array[15121] = 16'hdfc5;
mem_array[15120] = 16'h3c93;
mem_array[15123] = 16'h44a2;
mem_array[15122] = 16'h3d97;
mem_array[15125] = 16'h8153;
mem_array[15124] = 16'hbd0b;
mem_array[15127] = 16'h9911;
mem_array[15126] = 16'h3d6f;
mem_array[15129] = 16'h80a5;
mem_array[15128] = 16'h3db3;
mem_array[15131] = 16'h14b9;
mem_array[15130] = 16'hbd45;
mem_array[15133] = 16'h9efb;
mem_array[15132] = 16'h3dcb;
mem_array[15135] = 16'hde71;
mem_array[15134] = 16'hbc9b;
mem_array[15137] = 16'h157e;
mem_array[15136] = 16'h3d7a;
mem_array[15139] = 16'hd24a;
mem_array[15138] = 16'h3a18;
mem_array[15141] = 16'ha385;
mem_array[15140] = 16'hbcd2;
mem_array[15143] = 16'h3340;
mem_array[15142] = 16'hbd79;
mem_array[15145] = 16'he82e;
mem_array[15144] = 16'h3dbf;
mem_array[15147] = 16'hfbce;
mem_array[15146] = 16'hbce3;
mem_array[15149] = 16'hb02f;
mem_array[15148] = 16'hbc41;
mem_array[15151] = 16'hdc11;
mem_array[15150] = 16'hbe2d;
mem_array[15153] = 16'h663a;
mem_array[15152] = 16'h3c03;
mem_array[15155] = 16'he50d;
mem_array[15154] = 16'hbc88;
mem_array[15157] = 16'h9511;
mem_array[15156] = 16'h3e0e;
mem_array[15159] = 16'hc91f;
mem_array[15158] = 16'h3da1;
mem_array[15161] = 16'he471;
mem_array[15160] = 16'hbdfd;
mem_array[15163] = 16'hab18;
mem_array[15162] = 16'hbda4;
mem_array[15165] = 16'h20e1;
mem_array[15164] = 16'h3d4e;
mem_array[15167] = 16'h4417;
mem_array[15166] = 16'hbd7f;
mem_array[15169] = 16'h7b30;
mem_array[15168] = 16'h3b2f;
mem_array[15171] = 16'h3d48;
mem_array[15170] = 16'h3d39;
mem_array[15173] = 16'hd204;
mem_array[15172] = 16'hbd7c;
mem_array[15175] = 16'h88bf;
mem_array[15174] = 16'h3e19;
mem_array[15177] = 16'h166e;
mem_array[15176] = 16'h3c45;
mem_array[15179] = 16'h211e;
mem_array[15178] = 16'hbdf0;
mem_array[15181] = 16'h64ee;
mem_array[15180] = 16'h3d2d;
mem_array[15183] = 16'haf82;
mem_array[15182] = 16'h3fb9;
mem_array[15185] = 16'h2d71;
mem_array[15184] = 16'h3eea;
mem_array[15187] = 16'h3cf8;
mem_array[15186] = 16'h3d6c;
mem_array[15189] = 16'ha5bc;
mem_array[15188] = 16'h3e01;
mem_array[15191] = 16'h469e;
mem_array[15190] = 16'h3d31;
mem_array[15193] = 16'h99bf;
mem_array[15192] = 16'h3f49;
mem_array[15195] = 16'h0b75;
mem_array[15194] = 16'h3f66;
mem_array[15197] = 16'he8a7;
mem_array[15196] = 16'hbe8b;
mem_array[15199] = 16'h919d;
mem_array[15198] = 16'h3d8c;
mem_array[15201] = 16'hdfc5;
mem_array[15200] = 16'h3d7d;
mem_array[15203] = 16'hfec9;
mem_array[15202] = 16'h3db7;
mem_array[15205] = 16'hc1d8;
mem_array[15204] = 16'hbd11;
mem_array[15207] = 16'h66ad;
mem_array[15206] = 16'hbd8a;
mem_array[15209] = 16'hffd2;
mem_array[15208] = 16'hbe04;
mem_array[15211] = 16'h94b5;
mem_array[15210] = 16'h3d79;
mem_array[15213] = 16'h4879;
mem_array[15212] = 16'h3d58;
mem_array[15215] = 16'ha81a;
mem_array[15214] = 16'hbe5e;
mem_array[15217] = 16'h7854;
mem_array[15216] = 16'h3f40;
mem_array[15219] = 16'h7806;
mem_array[15218] = 16'h3e6b;
mem_array[15221] = 16'h9625;
mem_array[15220] = 16'hbf9b;
mem_array[15223] = 16'hcd0b;
mem_array[15222] = 16'h3e9a;
mem_array[15225] = 16'h43ff;
mem_array[15224] = 16'hbc2d;
mem_array[15227] = 16'h6a41;
mem_array[15226] = 16'hbf9c;
mem_array[15229] = 16'hbb01;
mem_array[15228] = 16'hbe5d;
mem_array[15231] = 16'h805e;
mem_array[15230] = 16'h3f7f;
mem_array[15233] = 16'h243b;
mem_array[15232] = 16'hbdd4;
mem_array[15235] = 16'hae69;
mem_array[15234] = 16'h3f24;
mem_array[15237] = 16'hef2f;
mem_array[15236] = 16'h3b00;
mem_array[15239] = 16'h4b5f;
mem_array[15238] = 16'hbfc2;
mem_array[15241] = 16'h0c8a;
mem_array[15240] = 16'h3f11;
mem_array[15243] = 16'h3d95;
mem_array[15242] = 16'hbf04;
mem_array[15245] = 16'h488d;
mem_array[15244] = 16'h3e87;
mem_array[15247] = 16'h07c5;
mem_array[15246] = 16'h3ec2;
mem_array[15249] = 16'h57fa;
mem_array[15248] = 16'h3d30;
mem_array[15251] = 16'hb24f;
mem_array[15250] = 16'h3ba6;
mem_array[15253] = 16'h65f2;
mem_array[15252] = 16'hbf05;
mem_array[15255] = 16'heb62;
mem_array[15254] = 16'hbf0a;
mem_array[15257] = 16'hd4aa;
mem_array[15256] = 16'hbef8;
mem_array[15259] = 16'he148;
mem_array[15258] = 16'h3e35;
mem_array[15261] = 16'h86a9;
mem_array[15260] = 16'hbda9;
mem_array[15263] = 16'hde94;
mem_array[15262] = 16'hbb32;
mem_array[15265] = 16'hb490;
mem_array[15264] = 16'h3ea4;
mem_array[15267] = 16'h457b;
mem_array[15266] = 16'hbf8e;
mem_array[15269] = 16'h7a97;
mem_array[15268] = 16'h3d84;
mem_array[15271] = 16'hdd15;
mem_array[15270] = 16'hbf37;
mem_array[15273] = 16'h0f84;
mem_array[15272] = 16'hbea4;
mem_array[15275] = 16'h1b75;
mem_array[15274] = 16'h3d61;
mem_array[15277] = 16'h962e;
mem_array[15276] = 16'h3cad;
mem_array[15279] = 16'hdbe3;
mem_array[15278] = 16'h3eea;
mem_array[15281] = 16'hf911;
mem_array[15280] = 16'h3ec6;
mem_array[15283] = 16'h9541;
mem_array[15282] = 16'h3f39;
mem_array[15285] = 16'hc01c;
mem_array[15284] = 16'h3d96;
mem_array[15287] = 16'hfa55;
mem_array[15286] = 16'h3f06;
mem_array[15289] = 16'h7040;
mem_array[15288] = 16'h3cf2;
mem_array[15291] = 16'h7dfa;
mem_array[15290] = 16'h3df3;
mem_array[15293] = 16'h72ae;
mem_array[15292] = 16'hbe6c;
mem_array[15295] = 16'haf09;
mem_array[15294] = 16'hbc22;
mem_array[15297] = 16'h0067;
mem_array[15296] = 16'hbe99;
mem_array[15299] = 16'h1d7f;
mem_array[15298] = 16'h3b5b;
mem_array[15301] = 16'h237b;
mem_array[15300] = 16'h3f42;
mem_array[15303] = 16'hd571;
mem_array[15302] = 16'hbd9f;
mem_array[15305] = 16'hb41b;
mem_array[15304] = 16'hbe95;
mem_array[15307] = 16'h3fcc;
mem_array[15306] = 16'hbf7e;
mem_array[15309] = 16'hbbbe;
mem_array[15308] = 16'h3ee4;
mem_array[15311] = 16'hde79;
mem_array[15310] = 16'hbee2;
mem_array[15313] = 16'h7398;
mem_array[15312] = 16'h3f1c;
mem_array[15315] = 16'h8f26;
mem_array[15314] = 16'h3e96;
mem_array[15317] = 16'h15b4;
mem_array[15316] = 16'h3eb1;
mem_array[15319] = 16'heb9e;
mem_array[15318] = 16'hbf17;
mem_array[15321] = 16'h07c7;
mem_array[15320] = 16'h3c0c;
mem_array[15323] = 16'hbe71;
mem_array[15322] = 16'h3be6;
mem_array[15325] = 16'h486b;
mem_array[15324] = 16'h3f15;
mem_array[15327] = 16'h2db9;
mem_array[15326] = 16'hbe67;
mem_array[15329] = 16'h922a;
mem_array[15328] = 16'h3e95;
mem_array[15331] = 16'h3c20;
mem_array[15330] = 16'hbed7;
mem_array[15333] = 16'h9b2c;
mem_array[15332] = 16'h3f6c;
mem_array[15335] = 16'heff5;
mem_array[15334] = 16'hbe2d;
mem_array[15337] = 16'h309d;
mem_array[15336] = 16'h3e75;
mem_array[15339] = 16'h2257;
mem_array[15338] = 16'hbe68;
mem_array[15341] = 16'he4e5;
mem_array[15340] = 16'hbf9b;
mem_array[15343] = 16'h4ab6;
mem_array[15342] = 16'h3e93;
mem_array[15345] = 16'hb866;
mem_array[15344] = 16'h3e21;
mem_array[15347] = 16'h802c;
mem_array[15346] = 16'hbd0b;
mem_array[15349] = 16'h9e4b;
mem_array[15348] = 16'h3f27;
mem_array[15351] = 16'hbe33;
mem_array[15350] = 16'h3ec1;
mem_array[15353] = 16'hf4a3;
mem_array[15352] = 16'h3eda;
mem_array[15355] = 16'he533;
mem_array[15354] = 16'h3d80;
mem_array[15357] = 16'h543b;
mem_array[15356] = 16'hbdb0;
mem_array[15359] = 16'he96f;
mem_array[15358] = 16'hbfa4;
mem_array[15361] = 16'h0b5c;
mem_array[15360] = 16'h3eef;
mem_array[15363] = 16'hcea4;
mem_array[15362] = 16'h3e92;
mem_array[15365] = 16'hacf3;
mem_array[15364] = 16'h3dce;
mem_array[15367] = 16'hd749;
mem_array[15366] = 16'hbd00;
mem_array[15369] = 16'h4eed;
mem_array[15368] = 16'hbf5b;
mem_array[15371] = 16'h76ff;
mem_array[15370] = 16'hbf4c;
mem_array[15373] = 16'h9dd0;
mem_array[15372] = 16'h3f34;
mem_array[15375] = 16'hccf2;
mem_array[15374] = 16'hbe28;
mem_array[15377] = 16'h7f68;
mem_array[15376] = 16'hbf05;
mem_array[15379] = 16'h3baa;
mem_array[15378] = 16'hbdbc;
mem_array[15381] = 16'h002c;
mem_array[15380] = 16'hbd18;
mem_array[15383] = 16'h9c0c;
mem_array[15382] = 16'h3d1e;
mem_array[15385] = 16'hee12;
mem_array[15384] = 16'hbefc;
mem_array[15387] = 16'h2d34;
mem_array[15386] = 16'h3f13;
mem_array[15389] = 16'ha185;
mem_array[15388] = 16'h3e1b;
mem_array[15391] = 16'hacbc;
mem_array[15390] = 16'hbe45;
mem_array[15393] = 16'h6f9b;
mem_array[15392] = 16'h3e59;
mem_array[15395] = 16'haad2;
mem_array[15394] = 16'hbe33;
mem_array[15397] = 16'h5632;
mem_array[15396] = 16'h3e6c;
mem_array[15399] = 16'h7da2;
mem_array[15398] = 16'hbed0;
mem_array[15401] = 16'h8536;
mem_array[15400] = 16'hbe38;
mem_array[15403] = 16'h2e63;
mem_array[15402] = 16'hbde2;
mem_array[15405] = 16'he4af;
mem_array[15404] = 16'hbc60;
mem_array[15407] = 16'h2439;
mem_array[15406] = 16'h3d5d;
mem_array[15409] = 16'hce14;
mem_array[15408] = 16'h3e39;
mem_array[15411] = 16'h2f3d;
mem_array[15410] = 16'h3ea7;
mem_array[15413] = 16'h3972;
mem_array[15412] = 16'hbe55;
mem_array[15415] = 16'h59ec;
mem_array[15414] = 16'h3d91;
mem_array[15417] = 16'h5022;
mem_array[15416] = 16'hbefd;
mem_array[15419] = 16'h0bc6;
mem_array[15418] = 16'hbf15;
mem_array[15421] = 16'hd64e;
mem_array[15420] = 16'h3e7f;
mem_array[15423] = 16'hba18;
mem_array[15422] = 16'h3ebf;
mem_array[15425] = 16'h9112;
mem_array[15424] = 16'h3ec1;
mem_array[15427] = 16'h15ee;
mem_array[15426] = 16'hbe3e;
mem_array[15429] = 16'h7fa6;
mem_array[15428] = 16'hbe45;
mem_array[15431] = 16'hffad;
mem_array[15430] = 16'hbe01;
mem_array[15433] = 16'hb6b2;
mem_array[15432] = 16'h3f22;
mem_array[15435] = 16'hec50;
mem_array[15434] = 16'hbd9f;
mem_array[15437] = 16'h7f04;
mem_array[15436] = 16'h3e34;
mem_array[15439] = 16'h46ce;
mem_array[15438] = 16'h3e5c;
mem_array[15441] = 16'hc16e;
mem_array[15440] = 16'hbd99;
mem_array[15443] = 16'h2255;
mem_array[15442] = 16'hbce3;
mem_array[15445] = 16'h738d;
mem_array[15444] = 16'hbec0;
mem_array[15447] = 16'h06d7;
mem_array[15446] = 16'hbe54;
mem_array[15449] = 16'hb915;
mem_array[15448] = 16'hbec6;
mem_array[15451] = 16'h6fa8;
mem_array[15450] = 16'h3e45;
mem_array[15453] = 16'h8aff;
mem_array[15452] = 16'hbe5a;
mem_array[15455] = 16'hd7ad;
mem_array[15454] = 16'h3ed0;
mem_array[15457] = 16'hb3d7;
mem_array[15456] = 16'hbe58;
mem_array[15459] = 16'h7aeb;
mem_array[15458] = 16'hbc90;
mem_array[15461] = 16'hd550;
mem_array[15460] = 16'hbf2f;
mem_array[15463] = 16'ha024;
mem_array[15462] = 16'hbddc;
mem_array[15465] = 16'haa66;
mem_array[15464] = 16'hbf26;
mem_array[15467] = 16'h3267;
mem_array[15466] = 16'hbd4e;
mem_array[15469] = 16'h4fec;
mem_array[15468] = 16'hbd3f;
mem_array[15471] = 16'h4e0f;
mem_array[15470] = 16'hbda2;
mem_array[15473] = 16'hc506;
mem_array[15472] = 16'hbdf2;
mem_array[15475] = 16'hba32;
mem_array[15474] = 16'hbf42;
mem_array[15477] = 16'h9617;
mem_array[15476] = 16'h3dcd;
mem_array[15479] = 16'hf1fc;
mem_array[15478] = 16'h3e01;
mem_array[15481] = 16'h4f2c;
mem_array[15480] = 16'h3f17;
mem_array[15483] = 16'he5ac;
mem_array[15482] = 16'h3e86;
mem_array[15485] = 16'hc01f;
mem_array[15484] = 16'h3c16;
mem_array[15487] = 16'h74b7;
mem_array[15486] = 16'hbd30;
mem_array[15489] = 16'h979e;
mem_array[15488] = 16'h3c76;
mem_array[15491] = 16'hd6de;
mem_array[15490] = 16'h3efa;
mem_array[15493] = 16'h61d0;
mem_array[15492] = 16'h3e55;
mem_array[15495] = 16'hb317;
mem_array[15494] = 16'h3e97;
mem_array[15497] = 16'h9bed;
mem_array[15496] = 16'hbe70;
mem_array[15499] = 16'h9336;
mem_array[15498] = 16'h3ee3;
mem_array[15501] = 16'hc41a;
mem_array[15500] = 16'hbd8b;
mem_array[15503] = 16'haf3f;
mem_array[15502] = 16'hbb94;
mem_array[15505] = 16'h27ef;
mem_array[15504] = 16'h3b94;
mem_array[15507] = 16'h82fe;
mem_array[15506] = 16'hbf2a;
mem_array[15509] = 16'h28f6;
mem_array[15508] = 16'hbcfa;
mem_array[15511] = 16'h34b0;
mem_array[15510] = 16'h3e20;
mem_array[15513] = 16'h2b38;
mem_array[15512] = 16'hbeef;
mem_array[15515] = 16'h050b;
mem_array[15514] = 16'hbe36;
mem_array[15517] = 16'h4c87;
mem_array[15516] = 16'h3ecb;
mem_array[15519] = 16'h4e6e;
mem_array[15518] = 16'hbe31;
mem_array[15521] = 16'h9cc6;
mem_array[15520] = 16'hbe9d;
mem_array[15523] = 16'hd6c2;
mem_array[15522] = 16'h3ea8;
mem_array[15525] = 16'h71d1;
mem_array[15524] = 16'hbf4d;
mem_array[15527] = 16'hab9a;
mem_array[15526] = 16'h3d4c;
mem_array[15529] = 16'h4a1c;
mem_array[15528] = 16'h3d29;
mem_array[15531] = 16'hfc2d;
mem_array[15530] = 16'h3f0a;
mem_array[15533] = 16'hb7ad;
mem_array[15532] = 16'h3d96;
mem_array[15535] = 16'h5d6a;
mem_array[15534] = 16'hbe48;
mem_array[15537] = 16'h8323;
mem_array[15536] = 16'h3e26;
mem_array[15539] = 16'h9443;
mem_array[15538] = 16'h3e50;
mem_array[15541] = 16'hfde8;
mem_array[15540] = 16'h3f13;
mem_array[15543] = 16'h3483;
mem_array[15542] = 16'h3e91;
mem_array[15545] = 16'h453a;
mem_array[15544] = 16'hbded;
mem_array[15547] = 16'h696a;
mem_array[15546] = 16'hbe8b;
mem_array[15549] = 16'h563b;
mem_array[15548] = 16'h3eae;
mem_array[15551] = 16'hb487;
mem_array[15550] = 16'hbedf;
mem_array[15553] = 16'h08a5;
mem_array[15552] = 16'hbc13;
mem_array[15555] = 16'h4484;
mem_array[15554] = 16'hbef8;
mem_array[15557] = 16'h420b;
mem_array[15556] = 16'h3d57;
mem_array[15559] = 16'h815a;
mem_array[15558] = 16'h3e22;
mem_array[15561] = 16'h87b2;
mem_array[15560] = 16'h3c86;
mem_array[15563] = 16'h807a;
mem_array[15562] = 16'hbddd;
mem_array[15565] = 16'h2578;
mem_array[15564] = 16'hbe09;
mem_array[15567] = 16'h2899;
mem_array[15566] = 16'hbe9d;
mem_array[15569] = 16'he168;
mem_array[15568] = 16'h3de3;
mem_array[15571] = 16'h7378;
mem_array[15570] = 16'h3deb;
mem_array[15573] = 16'h0bda;
mem_array[15572] = 16'h3e03;
mem_array[15575] = 16'h00eb;
mem_array[15574] = 16'hbdcf;
mem_array[15577] = 16'h77a6;
mem_array[15576] = 16'h3e02;
mem_array[15579] = 16'hb2cd;
mem_array[15578] = 16'hbe72;
mem_array[15581] = 16'h8d83;
mem_array[15580] = 16'h3e0d;
mem_array[15583] = 16'h0ec0;
mem_array[15582] = 16'h3ddf;
mem_array[15585] = 16'h483a;
mem_array[15584] = 16'h3ded;
mem_array[15587] = 16'hd708;
mem_array[15586] = 16'h3dbd;
mem_array[15589] = 16'haf8e;
mem_array[15588] = 16'h3e8d;
mem_array[15591] = 16'h2786;
mem_array[15590] = 16'h3f0c;
mem_array[15593] = 16'h335d;
mem_array[15592] = 16'h3d79;
mem_array[15595] = 16'ha7de;
mem_array[15594] = 16'hbe9b;
mem_array[15597] = 16'h0635;
mem_array[15596] = 16'hbd3e;
mem_array[15599] = 16'h1ace;
mem_array[15598] = 16'hbe79;
mem_array[15601] = 16'hc2dd;
mem_array[15600] = 16'h3eac;
mem_array[15603] = 16'h32d3;
mem_array[15602] = 16'h3d26;
mem_array[15605] = 16'h231b;
mem_array[15604] = 16'hbdce;
mem_array[15607] = 16'h9dfb;
mem_array[15606] = 16'hbecf;
mem_array[15609] = 16'h658f;
mem_array[15608] = 16'h3d08;
mem_array[15611] = 16'hd27e;
mem_array[15610] = 16'hbecb;
mem_array[15613] = 16'h1b51;
mem_array[15612] = 16'h3d83;
mem_array[15615] = 16'hc987;
mem_array[15614] = 16'hbf41;
mem_array[15617] = 16'h161d;
mem_array[15616] = 16'h3dd4;
mem_array[15619] = 16'h28e0;
mem_array[15618] = 16'hbb8f;
mem_array[15621] = 16'h13c6;
mem_array[15620] = 16'hbc92;
mem_array[15623] = 16'h8fb0;
mem_array[15622] = 16'h3ceb;
mem_array[15625] = 16'h1e50;
mem_array[15624] = 16'hbd28;
mem_array[15627] = 16'h9549;
mem_array[15626] = 16'hbe93;
mem_array[15629] = 16'h6740;
mem_array[15628] = 16'h3e7d;
mem_array[15631] = 16'hebfb;
mem_array[15630] = 16'h3e31;
mem_array[15633] = 16'hbd9a;
mem_array[15632] = 16'hbdcf;
mem_array[15635] = 16'h9c4b;
mem_array[15634] = 16'h3e80;
mem_array[15637] = 16'hafc6;
mem_array[15636] = 16'hbe08;
mem_array[15639] = 16'h217f;
mem_array[15638] = 16'hbcf3;
mem_array[15641] = 16'haee0;
mem_array[15640] = 16'h3c5b;
mem_array[15643] = 16'h714c;
mem_array[15642] = 16'h3eca;
mem_array[15645] = 16'h44ca;
mem_array[15644] = 16'h3e87;
mem_array[15647] = 16'h272c;
mem_array[15646] = 16'hbd5d;
mem_array[15649] = 16'h1058;
mem_array[15648] = 16'h3e82;
mem_array[15651] = 16'hcf54;
mem_array[15650] = 16'h3d1a;
mem_array[15653] = 16'hf048;
mem_array[15652] = 16'h3d3f;
mem_array[15655] = 16'hd27a;
mem_array[15654] = 16'hbd32;
mem_array[15657] = 16'hf883;
mem_array[15656] = 16'h3e4b;
mem_array[15659] = 16'h172c;
mem_array[15658] = 16'hbdbb;
mem_array[15661] = 16'h62f6;
mem_array[15660] = 16'h3eca;
mem_array[15663] = 16'hc12d;
mem_array[15662] = 16'h3dfc;
mem_array[15665] = 16'hb5f8;
mem_array[15664] = 16'h3e81;
mem_array[15667] = 16'hce66;
mem_array[15666] = 16'hbe13;
mem_array[15669] = 16'hb122;
mem_array[15668] = 16'hbdbf;
mem_array[15671] = 16'hc398;
mem_array[15670] = 16'h3e14;
mem_array[15673] = 16'h3120;
mem_array[15672] = 16'hbef6;
mem_array[15675] = 16'hfecd;
mem_array[15674] = 16'hbf67;
mem_array[15677] = 16'h3180;
mem_array[15676] = 16'h3e5c;
mem_array[15679] = 16'hfb9a;
mem_array[15678] = 16'hbe32;
mem_array[15681] = 16'h42f5;
mem_array[15680] = 16'hbda1;
mem_array[15683] = 16'ha827;
mem_array[15682] = 16'hbdb7;
mem_array[15685] = 16'hee10;
mem_array[15684] = 16'hbe7f;
mem_array[15687] = 16'h4490;
mem_array[15686] = 16'hbdcf;
mem_array[15689] = 16'h0462;
mem_array[15688] = 16'hbeab;
mem_array[15691] = 16'ha135;
mem_array[15690] = 16'h3e03;
mem_array[15693] = 16'h4f3c;
mem_array[15692] = 16'h3d50;
mem_array[15695] = 16'h3b04;
mem_array[15694] = 16'h3d90;
mem_array[15697] = 16'h959f;
mem_array[15696] = 16'h3cdc;
mem_array[15699] = 16'h13c2;
mem_array[15698] = 16'h3dc1;
mem_array[15701] = 16'hfb2c;
mem_array[15700] = 16'hbee2;
mem_array[15703] = 16'h9c76;
mem_array[15702] = 16'h3d1d;
mem_array[15705] = 16'h6b1e;
mem_array[15704] = 16'hbea6;
mem_array[15707] = 16'h5a64;
mem_array[15706] = 16'hbe20;
mem_array[15709] = 16'h5381;
mem_array[15708] = 16'h3e41;
mem_array[15711] = 16'h9d59;
mem_array[15710] = 16'h3ed3;
mem_array[15713] = 16'h4851;
mem_array[15712] = 16'h3d49;
mem_array[15715] = 16'h8fbb;
mem_array[15714] = 16'hbe16;
mem_array[15717] = 16'hc1fd;
mem_array[15716] = 16'hbc98;
mem_array[15719] = 16'h4665;
mem_array[15718] = 16'hbd98;
mem_array[15721] = 16'h5c75;
mem_array[15720] = 16'h3ef3;
mem_array[15723] = 16'h1d39;
mem_array[15722] = 16'hbe96;
mem_array[15725] = 16'hd43d;
mem_array[15724] = 16'h3e81;
mem_array[15727] = 16'h8452;
mem_array[15726] = 16'h3b95;
mem_array[15729] = 16'h9db7;
mem_array[15728] = 16'hbda5;
mem_array[15731] = 16'h15c5;
mem_array[15730] = 16'hbdb1;
mem_array[15733] = 16'h0a6a;
mem_array[15732] = 16'hbf80;
mem_array[15735] = 16'h366c;
mem_array[15734] = 16'hbf16;
mem_array[15737] = 16'hf9fb;
mem_array[15736] = 16'h3d08;
mem_array[15739] = 16'h2b72;
mem_array[15738] = 16'hbe28;
mem_array[15741] = 16'hd976;
mem_array[15740] = 16'hbdff;
mem_array[15743] = 16'h8760;
mem_array[15742] = 16'hbdef;
mem_array[15745] = 16'ha973;
mem_array[15744] = 16'hbe48;
mem_array[15747] = 16'hd396;
mem_array[15746] = 16'hbec2;
mem_array[15749] = 16'hce3c;
mem_array[15748] = 16'hbea0;
mem_array[15751] = 16'hbdf9;
mem_array[15750] = 16'h3e58;
mem_array[15753] = 16'h2285;
mem_array[15752] = 16'hbeca;
mem_array[15755] = 16'hae0e;
mem_array[15754] = 16'hbd1d;
mem_array[15757] = 16'hf83c;
mem_array[15756] = 16'h3d8c;
mem_array[15759] = 16'h009e;
mem_array[15758] = 16'hbe67;
mem_array[15761] = 16'h1af6;
mem_array[15760] = 16'hbda7;
mem_array[15763] = 16'h9c9a;
mem_array[15762] = 16'h3e26;
mem_array[15765] = 16'h332c;
mem_array[15764] = 16'h3cee;
mem_array[15767] = 16'he78b;
mem_array[15766] = 16'h3de8;
mem_array[15769] = 16'h13ad;
mem_array[15768] = 16'h3d91;
mem_array[15771] = 16'h852b;
mem_array[15770] = 16'h3e81;
mem_array[15773] = 16'h720c;
mem_array[15772] = 16'h3de1;
mem_array[15775] = 16'h6b50;
mem_array[15774] = 16'hbe07;
mem_array[15777] = 16'h890d;
mem_array[15776] = 16'hbd15;
mem_array[15779] = 16'hd4e0;
mem_array[15778] = 16'hbf1b;
mem_array[15781] = 16'hef1d;
mem_array[15780] = 16'hbece;
mem_array[15783] = 16'h1728;
mem_array[15782] = 16'h3d93;
mem_array[15785] = 16'h99a1;
mem_array[15784] = 16'h3e67;
mem_array[15787] = 16'h2078;
mem_array[15786] = 16'hbea2;
mem_array[15789] = 16'h5a02;
mem_array[15788] = 16'hbdee;
mem_array[15791] = 16'h3cf1;
mem_array[15790] = 16'h3e87;
mem_array[15793] = 16'h8308;
mem_array[15792] = 16'hbf4b;
mem_array[15795] = 16'h7dfa;
mem_array[15794] = 16'hbe93;
mem_array[15797] = 16'h3bf3;
mem_array[15796] = 16'h3e49;
mem_array[15799] = 16'h8dd8;
mem_array[15798] = 16'hbec5;
mem_array[15801] = 16'hbb15;
mem_array[15800] = 16'h3cec;
mem_array[15803] = 16'h2fdb;
mem_array[15802] = 16'h38ce;
mem_array[15805] = 16'h7dfd;
mem_array[15804] = 16'hbea0;
mem_array[15807] = 16'h3828;
mem_array[15806] = 16'h3e8b;
mem_array[15809] = 16'ha6b4;
mem_array[15808] = 16'hbe2a;
mem_array[15811] = 16'hf55b;
mem_array[15810] = 16'hbd14;
mem_array[15813] = 16'h09fe;
mem_array[15812] = 16'hbe94;
mem_array[15815] = 16'h222f;
mem_array[15814] = 16'h3ea3;
mem_array[15817] = 16'he769;
mem_array[15816] = 16'h3c93;
mem_array[15819] = 16'hab14;
mem_array[15818] = 16'hbedf;
mem_array[15821] = 16'hd714;
mem_array[15820] = 16'hbdd0;
mem_array[15823] = 16'h01bd;
mem_array[15822] = 16'h3d9b;
mem_array[15825] = 16'h6927;
mem_array[15824] = 16'hbf1c;
mem_array[15827] = 16'h998b;
mem_array[15826] = 16'hbcb1;
mem_array[15829] = 16'hb477;
mem_array[15828] = 16'h3ecf;
mem_array[15831] = 16'hb76f;
mem_array[15830] = 16'h3e82;
mem_array[15833] = 16'hc65e;
mem_array[15832] = 16'h3e13;
mem_array[15835] = 16'h8fd3;
mem_array[15834] = 16'h3c4d;
mem_array[15837] = 16'hc33e;
mem_array[15836] = 16'h3e66;
mem_array[15839] = 16'h97a5;
mem_array[15838] = 16'hbed8;
mem_array[15841] = 16'h02e4;
mem_array[15840] = 16'hbef9;
mem_array[15843] = 16'h62a6;
mem_array[15842] = 16'h3d4f;
mem_array[15845] = 16'ha918;
mem_array[15844] = 16'h3eb5;
mem_array[15847] = 16'hec58;
mem_array[15846] = 16'hbde1;
mem_array[15849] = 16'hb7cb;
mem_array[15848] = 16'hbda8;
mem_array[15851] = 16'hfd9c;
mem_array[15850] = 16'hbcd4;
mem_array[15853] = 16'hfb02;
mem_array[15852] = 16'hbf3c;
mem_array[15855] = 16'h4a5f;
mem_array[15854] = 16'hbed3;
mem_array[15857] = 16'he313;
mem_array[15856] = 16'h3e17;
mem_array[15859] = 16'h1eb7;
mem_array[15858] = 16'hbdbc;
mem_array[15861] = 16'hbf14;
mem_array[15860] = 16'hbd6e;
mem_array[15863] = 16'h592b;
mem_array[15862] = 16'h3cf4;
mem_array[15865] = 16'h73dd;
mem_array[15864] = 16'hbe19;
mem_array[15867] = 16'h49ae;
mem_array[15866] = 16'h3cdb;
mem_array[15869] = 16'h1a04;
mem_array[15868] = 16'hbdbc;
mem_array[15871] = 16'h3f75;
mem_array[15870] = 16'h3e18;
mem_array[15873] = 16'h85a3;
mem_array[15872] = 16'hbc8b;
mem_array[15875] = 16'hc6a5;
mem_array[15874] = 16'h3e90;
mem_array[15877] = 16'h7106;
mem_array[15876] = 16'h3e8a;
mem_array[15879] = 16'h2815;
mem_array[15878] = 16'hbe32;
mem_array[15881] = 16'h1d93;
mem_array[15880] = 16'hbe90;
mem_array[15883] = 16'h8b3f;
mem_array[15882] = 16'h3e8b;
mem_array[15885] = 16'h48df;
mem_array[15884] = 16'hbdf2;
mem_array[15887] = 16'hed89;
mem_array[15886] = 16'h3e25;
mem_array[15889] = 16'h0084;
mem_array[15888] = 16'h3e9d;
mem_array[15891] = 16'h2441;
mem_array[15890] = 16'h3ef0;
mem_array[15893] = 16'h4e51;
mem_array[15892] = 16'hbdbc;
mem_array[15895] = 16'h1437;
mem_array[15894] = 16'h3e64;
mem_array[15897] = 16'h5a81;
mem_array[15896] = 16'h3ecc;
mem_array[15899] = 16'h2ff5;
mem_array[15898] = 16'hbeb2;
mem_array[15901] = 16'hcce9;
mem_array[15900] = 16'hbf61;
mem_array[15903] = 16'hae7b;
mem_array[15902] = 16'hbde0;
mem_array[15905] = 16'h8069;
mem_array[15904] = 16'h3c9a;
mem_array[15907] = 16'hf49f;
mem_array[15906] = 16'h3e43;
mem_array[15909] = 16'hf505;
mem_array[15908] = 16'hbe22;
mem_array[15911] = 16'hb990;
mem_array[15910] = 16'h3de7;
mem_array[15913] = 16'h0341;
mem_array[15912] = 16'hbe73;
mem_array[15915] = 16'h485f;
mem_array[15914] = 16'hbde6;
mem_array[15917] = 16'ha5dc;
mem_array[15916] = 16'h3e32;
mem_array[15919] = 16'h1df8;
mem_array[15918] = 16'h3ec3;
mem_array[15921] = 16'ha599;
mem_array[15920] = 16'hbd84;
mem_array[15923] = 16'h0383;
mem_array[15922] = 16'h3c1d;
mem_array[15925] = 16'hf06d;
mem_array[15924] = 16'hbdc0;
mem_array[15927] = 16'hb608;
mem_array[15926] = 16'hbea0;
mem_array[15929] = 16'hb8d7;
mem_array[15928] = 16'hbd93;
mem_array[15931] = 16'h4e91;
mem_array[15930] = 16'hbd2f;
mem_array[15933] = 16'h4a4b;
mem_array[15932] = 16'hbe17;
mem_array[15935] = 16'h1c8f;
mem_array[15934] = 16'h3db2;
mem_array[15937] = 16'h03d2;
mem_array[15936] = 16'hbbbe;
mem_array[15939] = 16'hb840;
mem_array[15938] = 16'h3dfe;
mem_array[15941] = 16'h9b38;
mem_array[15940] = 16'h3b40;
mem_array[15943] = 16'h5fb9;
mem_array[15942] = 16'h3c1a;
mem_array[15945] = 16'h4655;
mem_array[15944] = 16'hbdbf;
mem_array[15947] = 16'h1dc1;
mem_array[15946] = 16'h3d8b;
mem_array[15949] = 16'h5f14;
mem_array[15948] = 16'hbe3d;
mem_array[15951] = 16'hb62e;
mem_array[15950] = 16'h3ee8;
mem_array[15953] = 16'h89e3;
mem_array[15952] = 16'hbe9a;
mem_array[15955] = 16'h6fd3;
mem_array[15954] = 16'h3e22;
mem_array[15957] = 16'hc916;
mem_array[15956] = 16'h3c87;
mem_array[15959] = 16'h018f;
mem_array[15958] = 16'hbe7e;
mem_array[15961] = 16'h580a;
mem_array[15960] = 16'hbe93;
mem_array[15963] = 16'he4d9;
mem_array[15962] = 16'hbd2e;
mem_array[15965] = 16'h1a84;
mem_array[15964] = 16'hbe83;
mem_array[15967] = 16'h2fd2;
mem_array[15966] = 16'h3b8c;
mem_array[15969] = 16'hdd3c;
mem_array[15968] = 16'hbc78;
mem_array[15971] = 16'h88f4;
mem_array[15970] = 16'hbde9;
mem_array[15973] = 16'h1766;
mem_array[15972] = 16'h3c5c;
mem_array[15975] = 16'he22e;
mem_array[15974] = 16'hbdfa;
mem_array[15977] = 16'habfa;
mem_array[15976] = 16'h3f09;
mem_array[15979] = 16'h9e9e;
mem_array[15978] = 16'h3f32;
mem_array[15981] = 16'he63a;
mem_array[15980] = 16'h3d47;
mem_array[15983] = 16'h2ec0;
mem_array[15982] = 16'hbdbf;
mem_array[15985] = 16'h321f;
mem_array[15984] = 16'hbde1;
mem_array[15987] = 16'hd439;
mem_array[15986] = 16'hbe31;
mem_array[15989] = 16'h08b8;
mem_array[15988] = 16'hbd98;
mem_array[15991] = 16'h0580;
mem_array[15990] = 16'hbdf5;
mem_array[15993] = 16'hcefe;
mem_array[15992] = 16'hbbf6;
mem_array[15995] = 16'h1350;
mem_array[15994] = 16'hbffd;
mem_array[15997] = 16'hbf14;
mem_array[15996] = 16'h3e6f;
mem_array[15999] = 16'h524f;
mem_array[15998] = 16'hbf29;
mem_array[16001] = 16'h8449;
mem_array[16000] = 16'hbe0a;
mem_array[16003] = 16'h6433;
mem_array[16002] = 16'h3e5e;
mem_array[16005] = 16'hc265;
mem_array[16004] = 16'h3d24;
mem_array[16007] = 16'h160f;
mem_array[16006] = 16'hbd8b;
mem_array[16009] = 16'hb970;
mem_array[16008] = 16'hbe50;
mem_array[16011] = 16'hac07;
mem_array[16010] = 16'h3e4e;
mem_array[16013] = 16'h4a0a;
mem_array[16012] = 16'hbe2a;
mem_array[16015] = 16'ha81a;
mem_array[16014] = 16'h3aa1;
mem_array[16017] = 16'h497d;
mem_array[16016] = 16'hbd9b;
mem_array[16019] = 16'h4d45;
mem_array[16018] = 16'hbeab;
mem_array[16021] = 16'h465d;
mem_array[16020] = 16'h3e46;
mem_array[16023] = 16'h3dea;
mem_array[16022] = 16'hbe3d;
mem_array[16025] = 16'hc154;
mem_array[16024] = 16'hbe5a;
mem_array[16027] = 16'h3a3e;
mem_array[16026] = 16'h3da8;
mem_array[16029] = 16'h5157;
mem_array[16028] = 16'hbd84;
mem_array[16031] = 16'had57;
mem_array[16030] = 16'hbf3a;
mem_array[16033] = 16'h8497;
mem_array[16032] = 16'h3ecd;
mem_array[16035] = 16'hea6e;
mem_array[16034] = 16'hbd83;
mem_array[16037] = 16'h3f6a;
mem_array[16036] = 16'h3e6a;
mem_array[16039] = 16'hb257;
mem_array[16038] = 16'h3ea7;
mem_array[16041] = 16'hf983;
mem_array[16040] = 16'h3d26;
mem_array[16043] = 16'hef48;
mem_array[16042] = 16'hbda5;
mem_array[16045] = 16'h67cf;
mem_array[16044] = 16'hbdef;
mem_array[16047] = 16'hc17f;
mem_array[16046] = 16'hbe33;
mem_array[16049] = 16'h7acf;
mem_array[16048] = 16'hbe8a;
mem_array[16051] = 16'h7ab4;
mem_array[16050] = 16'hbb89;
mem_array[16053] = 16'h0a3f;
mem_array[16052] = 16'h3d70;
mem_array[16055] = 16'h867f;
mem_array[16054] = 16'hbdef;
mem_array[16057] = 16'hcf19;
mem_array[16056] = 16'h3e66;
mem_array[16059] = 16'ha596;
mem_array[16058] = 16'hbf03;
mem_array[16061] = 16'h845c;
mem_array[16060] = 16'h3e2a;
mem_array[16063] = 16'h3c89;
mem_array[16062] = 16'h3eef;
mem_array[16065] = 16'h3f78;
mem_array[16064] = 16'hbebd;
mem_array[16067] = 16'h661d;
mem_array[16066] = 16'hbda2;
mem_array[16069] = 16'h6012;
mem_array[16068] = 16'h3d06;
mem_array[16071] = 16'h62ac;
mem_array[16070] = 16'h3e44;
mem_array[16073] = 16'h8fe3;
mem_array[16072] = 16'hbe28;
mem_array[16075] = 16'hf715;
mem_array[16074] = 16'h3e7d;
mem_array[16077] = 16'h24da;
mem_array[16076] = 16'hbd95;
mem_array[16079] = 16'h9c7a;
mem_array[16078] = 16'h3e19;
mem_array[16081] = 16'hdb7a;
mem_array[16080] = 16'h3f24;
mem_array[16083] = 16'hb15b;
mem_array[16082] = 16'hbe1c;
mem_array[16085] = 16'h8754;
mem_array[16084] = 16'h3d0f;
mem_array[16087] = 16'h3135;
mem_array[16086] = 16'h3da6;
mem_array[16089] = 16'h0e9d;
mem_array[16088] = 16'h3c99;
mem_array[16091] = 16'h5e11;
mem_array[16090] = 16'hbf3b;
mem_array[16093] = 16'hf7bd;
mem_array[16092] = 16'h3e94;
mem_array[16095] = 16'h20e5;
mem_array[16094] = 16'h3de6;
mem_array[16097] = 16'h0244;
mem_array[16096] = 16'hbe04;
mem_array[16099] = 16'h796b;
mem_array[16098] = 16'h3dc5;
mem_array[16101] = 16'heb59;
mem_array[16100] = 16'hbcca;
mem_array[16103] = 16'h656d;
mem_array[16102] = 16'h3cef;
mem_array[16105] = 16'h0fcf;
mem_array[16104] = 16'h3e35;
mem_array[16107] = 16'h68d0;
mem_array[16106] = 16'h3dc3;
mem_array[16109] = 16'h85d6;
mem_array[16108] = 16'hbe8c;
mem_array[16111] = 16'hd82c;
mem_array[16110] = 16'h3e3e;
mem_array[16113] = 16'hb0a0;
mem_array[16112] = 16'h3f02;
mem_array[16115] = 16'h7b86;
mem_array[16114] = 16'h3ef9;
mem_array[16117] = 16'hf1f0;
mem_array[16116] = 16'hbd9c;
mem_array[16119] = 16'h7133;
mem_array[16118] = 16'hbdb3;
mem_array[16121] = 16'h8059;
mem_array[16120] = 16'hbe10;
mem_array[16123] = 16'hb743;
mem_array[16122] = 16'h3df2;
mem_array[16125] = 16'h1b22;
mem_array[16124] = 16'hbd9a;
mem_array[16127] = 16'hada2;
mem_array[16126] = 16'hbe05;
mem_array[16129] = 16'hdfb4;
mem_array[16128] = 16'h3d5d;
mem_array[16131] = 16'h3e10;
mem_array[16130] = 16'h3e0b;
mem_array[16133] = 16'h6b2f;
mem_array[16132] = 16'hbeb0;
mem_array[16135] = 16'h7348;
mem_array[16134] = 16'h3dff;
mem_array[16137] = 16'h6651;
mem_array[16136] = 16'hbde0;
mem_array[16139] = 16'h2ead;
mem_array[16138] = 16'hbd8a;
mem_array[16141] = 16'h6d8b;
mem_array[16140] = 16'h3dd5;
mem_array[16143] = 16'h758e;
mem_array[16142] = 16'h3dc2;
mem_array[16145] = 16'heedd;
mem_array[16144] = 16'h3e5a;
mem_array[16147] = 16'h3292;
mem_array[16146] = 16'h3dca;
mem_array[16149] = 16'h4641;
mem_array[16148] = 16'h3e3c;
mem_array[16151] = 16'h2e88;
mem_array[16150] = 16'hbefe;
mem_array[16153] = 16'h256e;
mem_array[16152] = 16'h3e67;
mem_array[16155] = 16'hdbbd;
mem_array[16154] = 16'hbd92;
mem_array[16157] = 16'hcd9b;
mem_array[16156] = 16'hbeb0;
mem_array[16159] = 16'h5fde;
mem_array[16158] = 16'hbec4;
mem_array[16161] = 16'h0989;
mem_array[16160] = 16'hbd88;
mem_array[16163] = 16'h8277;
mem_array[16162] = 16'h3d34;
mem_array[16165] = 16'hf9a8;
mem_array[16164] = 16'h3d91;
mem_array[16167] = 16'haa3b;
mem_array[16166] = 16'hbd8e;
mem_array[16169] = 16'h3434;
mem_array[16168] = 16'h3d15;
mem_array[16171] = 16'h9134;
mem_array[16170] = 16'h3e24;
mem_array[16173] = 16'hacf0;
mem_array[16172] = 16'hbe1b;
mem_array[16175] = 16'h86e1;
mem_array[16174] = 16'h3dec;
mem_array[16177] = 16'hd4e9;
mem_array[16176] = 16'h3e86;
mem_array[16179] = 16'h4a95;
mem_array[16178] = 16'hbddc;
mem_array[16181] = 16'h555a;
mem_array[16180] = 16'h3b2a;
mem_array[16183] = 16'hdc64;
mem_array[16182] = 16'h3e95;
mem_array[16185] = 16'h884c;
mem_array[16184] = 16'hbef4;
mem_array[16187] = 16'ha737;
mem_array[16186] = 16'hbe2b;
mem_array[16189] = 16'h4cfa;
mem_array[16188] = 16'h3e49;
mem_array[16191] = 16'h5c0b;
mem_array[16190] = 16'h3ed4;
mem_array[16193] = 16'h118b;
mem_array[16192] = 16'hbe7e;
mem_array[16195] = 16'hd7a1;
mem_array[16194] = 16'h3e8b;
mem_array[16197] = 16'h1d50;
mem_array[16196] = 16'hbeca;
mem_array[16199] = 16'h3a0c;
mem_array[16198] = 16'hbe71;
mem_array[16201] = 16'h1a49;
mem_array[16200] = 16'h3dc8;
mem_array[16203] = 16'h313a;
mem_array[16202] = 16'h3d4d;
mem_array[16205] = 16'h3e63;
mem_array[16204] = 16'hbe05;
mem_array[16207] = 16'h11ee;
mem_array[16206] = 16'h3e81;
mem_array[16209] = 16'hf23f;
mem_array[16208] = 16'h3c9c;
mem_array[16211] = 16'hc18b;
mem_array[16210] = 16'hbe02;
mem_array[16213] = 16'h54cb;
mem_array[16212] = 16'h3e41;
mem_array[16215] = 16'h4e3a;
mem_array[16214] = 16'h3d04;
mem_array[16217] = 16'h7a5e;
mem_array[16216] = 16'hbe5c;
mem_array[16219] = 16'hdc15;
mem_array[16218] = 16'hbe4b;
mem_array[16221] = 16'hc062;
mem_array[16220] = 16'hbc0a;
mem_array[16223] = 16'hbfab;
mem_array[16222] = 16'hbd02;
mem_array[16225] = 16'hdd04;
mem_array[16224] = 16'hbe82;
mem_array[16227] = 16'ha039;
mem_array[16226] = 16'h3e4b;
mem_array[16229] = 16'h2e46;
mem_array[16228] = 16'h3deb;
mem_array[16231] = 16'h787a;
mem_array[16230] = 16'h3e42;
mem_array[16233] = 16'h738c;
mem_array[16232] = 16'hbc91;
mem_array[16235] = 16'h7f6a;
mem_array[16234] = 16'hbe00;
mem_array[16237] = 16'hbe30;
mem_array[16236] = 16'hbdb0;
mem_array[16239] = 16'h7441;
mem_array[16238] = 16'h3d9b;
mem_array[16241] = 16'hd9b7;
mem_array[16240] = 16'hbe66;
mem_array[16243] = 16'hb0d5;
mem_array[16242] = 16'h3d34;
mem_array[16245] = 16'hb47b;
mem_array[16244] = 16'hbfe9;
mem_array[16247] = 16'h5fd7;
mem_array[16246] = 16'hbe01;
mem_array[16249] = 16'hf097;
mem_array[16248] = 16'h3d74;
mem_array[16251] = 16'h6b41;
mem_array[16250] = 16'h3e38;
mem_array[16253] = 16'h7873;
mem_array[16252] = 16'hbe92;
mem_array[16255] = 16'h6a21;
mem_array[16254] = 16'h3ef1;
mem_array[16257] = 16'h994f;
mem_array[16256] = 16'hbdc2;
mem_array[16259] = 16'h41d0;
mem_array[16258] = 16'hbec8;
mem_array[16261] = 16'h56c6;
mem_array[16260] = 16'hbe06;
mem_array[16263] = 16'hdf50;
mem_array[16262] = 16'hbdbf;
mem_array[16265] = 16'h23c1;
mem_array[16264] = 16'hbea4;
mem_array[16267] = 16'hd630;
mem_array[16266] = 16'h3f17;
mem_array[16269] = 16'h21e1;
mem_array[16268] = 16'h3e56;
mem_array[16271] = 16'h9315;
mem_array[16270] = 16'h3dd9;
mem_array[16273] = 16'hebe1;
mem_array[16272] = 16'h3e42;
mem_array[16275] = 16'h2db9;
mem_array[16274] = 16'hbdf2;
mem_array[16277] = 16'h1545;
mem_array[16276] = 16'hbe4f;
mem_array[16279] = 16'hea5e;
mem_array[16278] = 16'hbf04;
mem_array[16281] = 16'h1ea2;
mem_array[16280] = 16'hbcf0;
mem_array[16283] = 16'h7a41;
mem_array[16282] = 16'h3ccc;
mem_array[16285] = 16'h2bf8;
mem_array[16284] = 16'hbdc2;
mem_array[16287] = 16'h9c38;
mem_array[16286] = 16'h3c98;
mem_array[16289] = 16'h315d;
mem_array[16288] = 16'h3f0d;
mem_array[16291] = 16'h37cd;
mem_array[16290] = 16'h3e0c;
mem_array[16293] = 16'h43f7;
mem_array[16292] = 16'hbd46;
mem_array[16295] = 16'h53ca;
mem_array[16294] = 16'h3c8a;
mem_array[16297] = 16'he8ba;
mem_array[16296] = 16'hbd37;
mem_array[16299] = 16'hb069;
mem_array[16298] = 16'h3c04;
mem_array[16301] = 16'hbdd4;
mem_array[16300] = 16'h3d9b;
mem_array[16303] = 16'h2391;
mem_array[16302] = 16'hbbc7;
mem_array[16305] = 16'h4b40;
mem_array[16304] = 16'hc004;
mem_array[16307] = 16'h861f;
mem_array[16306] = 16'hbc5f;
mem_array[16309] = 16'h1eb3;
mem_array[16308] = 16'hbe22;
mem_array[16311] = 16'heffe;
mem_array[16310] = 16'h3d45;
mem_array[16313] = 16'hc928;
mem_array[16312] = 16'hbe1e;
mem_array[16315] = 16'h55ef;
mem_array[16314] = 16'h3dc7;
mem_array[16317] = 16'h933f;
mem_array[16316] = 16'h3dc2;
mem_array[16319] = 16'h6cad;
mem_array[16318] = 16'hbeaa;
mem_array[16321] = 16'he5f5;
mem_array[16320] = 16'hbec7;
mem_array[16323] = 16'hd640;
mem_array[16322] = 16'h3bf9;
mem_array[16325] = 16'hbf78;
mem_array[16324] = 16'hbe40;
mem_array[16327] = 16'hca55;
mem_array[16326] = 16'h3efb;
mem_array[16329] = 16'hb652;
mem_array[16328] = 16'h3e0b;
mem_array[16331] = 16'h72e9;
mem_array[16330] = 16'h3def;
mem_array[16333] = 16'hc7d6;
mem_array[16332] = 16'h3eb2;
mem_array[16335] = 16'h08b1;
mem_array[16334] = 16'hbd7b;
mem_array[16337] = 16'hd249;
mem_array[16336] = 16'h3e04;
mem_array[16339] = 16'h80ea;
mem_array[16338] = 16'hbfc2;
mem_array[16341] = 16'h2ab1;
mem_array[16340] = 16'h3cb4;
mem_array[16343] = 16'h3f0d;
mem_array[16342] = 16'hbcd5;
mem_array[16345] = 16'h0c57;
mem_array[16344] = 16'hbd68;
mem_array[16347] = 16'hd6ff;
mem_array[16346] = 16'hbe2d;
mem_array[16349] = 16'hf87a;
mem_array[16348] = 16'h3ea1;
mem_array[16351] = 16'h65fa;
mem_array[16350] = 16'hbda4;
mem_array[16353] = 16'h631e;
mem_array[16352] = 16'hbf02;
mem_array[16355] = 16'h8840;
mem_array[16354] = 16'h3e86;
mem_array[16357] = 16'haa83;
mem_array[16356] = 16'hbe81;
mem_array[16359] = 16'h94a4;
mem_array[16358] = 16'h3eb9;
mem_array[16361] = 16'hc1b0;
mem_array[16360] = 16'h3d3d;
mem_array[16363] = 16'h8a50;
mem_array[16362] = 16'hbe49;
mem_array[16365] = 16'h2c23;
mem_array[16364] = 16'hbfc4;
mem_array[16367] = 16'hf9c2;
mem_array[16366] = 16'h3d92;
mem_array[16369] = 16'hd657;
mem_array[16368] = 16'hbcee;
mem_array[16371] = 16'h2d1e;
mem_array[16370] = 16'h3e5f;
mem_array[16373] = 16'ha418;
mem_array[16372] = 16'hbec9;
mem_array[16375] = 16'h85e4;
mem_array[16374] = 16'h3992;
mem_array[16377] = 16'h9403;
mem_array[16376] = 16'hbcb8;
mem_array[16379] = 16'heb5c;
mem_array[16378] = 16'hbe93;
mem_array[16381] = 16'h42a3;
mem_array[16380] = 16'hbdb5;
mem_array[16383] = 16'h9a71;
mem_array[16382] = 16'h3ec6;
mem_array[16385] = 16'hcfea;
mem_array[16384] = 16'hbe6f;
mem_array[16387] = 16'h684f;
mem_array[16386] = 16'h3ca4;
mem_array[16389] = 16'h88fa;
mem_array[16388] = 16'h3d15;
mem_array[16391] = 16'hb866;
mem_array[16390] = 16'h3eb9;
mem_array[16393] = 16'hd118;
mem_array[16392] = 16'hbc58;
mem_array[16395] = 16'h5626;
mem_array[16394] = 16'hbd2f;
mem_array[16397] = 16'h1791;
mem_array[16396] = 16'hbe1e;
mem_array[16399] = 16'h7915;
mem_array[16398] = 16'h3eaa;
mem_array[16401] = 16'h0ae8;
mem_array[16400] = 16'h3cea;
mem_array[16403] = 16'h388f;
mem_array[16402] = 16'hbd69;
mem_array[16405] = 16'hb265;
mem_array[16404] = 16'hbe7d;
mem_array[16407] = 16'h661d;
mem_array[16406] = 16'hbdb3;
mem_array[16409] = 16'h0c9b;
mem_array[16408] = 16'h3ea0;
mem_array[16411] = 16'h8205;
mem_array[16410] = 16'h3e05;
mem_array[16413] = 16'h36bf;
mem_array[16412] = 16'h3d93;
mem_array[16415] = 16'h2c27;
mem_array[16414] = 16'h3d74;
mem_array[16417] = 16'hc799;
mem_array[16416] = 16'hbe10;
mem_array[16419] = 16'h2d5c;
mem_array[16418] = 16'h3e71;
mem_array[16421] = 16'h9097;
mem_array[16420] = 16'h3e19;
mem_array[16423] = 16'h4472;
mem_array[16422] = 16'h3d3a;
mem_array[16425] = 16'h995b;
mem_array[16424] = 16'hbfb6;
mem_array[16427] = 16'h17bc;
mem_array[16426] = 16'hbc8e;
mem_array[16429] = 16'hb4db;
mem_array[16428] = 16'hbe95;
mem_array[16431] = 16'h4a84;
mem_array[16430] = 16'h3eb6;
mem_array[16433] = 16'h7606;
mem_array[16432] = 16'hbeee;
mem_array[16435] = 16'h8e2d;
mem_array[16434] = 16'h3e29;
mem_array[16437] = 16'h7a63;
mem_array[16436] = 16'hbe73;
mem_array[16439] = 16'hcf3f;
mem_array[16438] = 16'hbf0a;
mem_array[16441] = 16'h971c;
mem_array[16440] = 16'h3e99;
mem_array[16443] = 16'hb3f7;
mem_array[16442] = 16'h3f00;
mem_array[16445] = 16'hff9b;
mem_array[16444] = 16'hbe1b;
mem_array[16447] = 16'h387a;
mem_array[16446] = 16'h3e20;
mem_array[16449] = 16'he259;
mem_array[16448] = 16'hbb97;
mem_array[16451] = 16'h376d;
mem_array[16450] = 16'h3f13;
mem_array[16453] = 16'hbf32;
mem_array[16452] = 16'hbd9c;
mem_array[16455] = 16'hf72b;
mem_array[16454] = 16'hbd97;
mem_array[16457] = 16'hd72b;
mem_array[16456] = 16'hbe5d;
mem_array[16459] = 16'h707f;
mem_array[16458] = 16'hbedd;
mem_array[16461] = 16'hff00;
mem_array[16460] = 16'hbd86;
mem_array[16463] = 16'h1078;
mem_array[16462] = 16'h3cc4;
mem_array[16465] = 16'he34e;
mem_array[16464] = 16'hbf02;
mem_array[16467] = 16'h4ebb;
mem_array[16466] = 16'h3d91;
mem_array[16469] = 16'hc68d;
mem_array[16468] = 16'hbdd7;
mem_array[16471] = 16'haa06;
mem_array[16470] = 16'h3ea4;
mem_array[16473] = 16'h32b4;
mem_array[16472] = 16'h3edc;
mem_array[16475] = 16'h0127;
mem_array[16474] = 16'h3e1f;
mem_array[16477] = 16'h64fd;
mem_array[16476] = 16'h3d8e;
mem_array[16479] = 16'h7026;
mem_array[16478] = 16'h3e80;
mem_array[16481] = 16'h7f70;
mem_array[16480] = 16'hba07;
mem_array[16483] = 16'hd34c;
mem_array[16482] = 16'h3d7c;
mem_array[16485] = 16'haaac;
mem_array[16484] = 16'hbf51;
mem_array[16487] = 16'h2869;
mem_array[16486] = 16'hba52;
mem_array[16489] = 16'h8662;
mem_array[16488] = 16'h3f24;
mem_array[16491] = 16'h8a27;
mem_array[16490] = 16'h3e1d;
mem_array[16493] = 16'hec2a;
mem_array[16492] = 16'h3daa;
mem_array[16495] = 16'h2e88;
mem_array[16494] = 16'h3f3e;
mem_array[16497] = 16'h6f24;
mem_array[16496] = 16'hbef6;
mem_array[16499] = 16'h1ee0;
mem_array[16498] = 16'hbfab;
mem_array[16501] = 16'h9a05;
mem_array[16500] = 16'hbea7;
mem_array[16503] = 16'h1f64;
mem_array[16502] = 16'h3e82;
mem_array[16505] = 16'h1bbc;
mem_array[16504] = 16'h3e39;
mem_array[16507] = 16'h5ce7;
mem_array[16506] = 16'h3ee3;
mem_array[16509] = 16'h6594;
mem_array[16508] = 16'hbea0;
mem_array[16511] = 16'h6fd0;
mem_array[16510] = 16'h3e74;
mem_array[16513] = 16'he092;
mem_array[16512] = 16'hbfd6;
mem_array[16515] = 16'hd3a9;
mem_array[16514] = 16'hbe86;
mem_array[16517] = 16'h2041;
mem_array[16516] = 16'hbd88;
mem_array[16519] = 16'h1989;
mem_array[16518] = 16'hbe2f;
mem_array[16521] = 16'h8fa5;
mem_array[16520] = 16'h3c90;
mem_array[16523] = 16'hdf7b;
mem_array[16522] = 16'h3b47;
mem_array[16525] = 16'he3d0;
mem_array[16524] = 16'hbe98;
mem_array[16527] = 16'h3bdc;
mem_array[16526] = 16'hbe12;
mem_array[16529] = 16'hd903;
mem_array[16528] = 16'h3efe;
mem_array[16531] = 16'hdd4b;
mem_array[16530] = 16'hbded;
mem_array[16533] = 16'hdfa5;
mem_array[16532] = 16'hbedb;
mem_array[16535] = 16'h6614;
mem_array[16534] = 16'hbcb6;
mem_array[16537] = 16'ha938;
mem_array[16536] = 16'hbe5c;
mem_array[16539] = 16'hf196;
mem_array[16538] = 16'h3d29;
mem_array[16541] = 16'h109b;
mem_array[16540] = 16'hbd7e;
mem_array[16543] = 16'hb578;
mem_array[16542] = 16'hbe26;
mem_array[16545] = 16'h4edf;
mem_array[16544] = 16'hbf4b;
mem_array[16547] = 16'hd809;
mem_array[16546] = 16'hbe4d;
mem_array[16549] = 16'h11d6;
mem_array[16548] = 16'h3eb4;
mem_array[16551] = 16'he810;
mem_array[16550] = 16'h3c04;
mem_array[16553] = 16'h09c0;
mem_array[16552] = 16'h3eba;
mem_array[16555] = 16'hf7de;
mem_array[16554] = 16'h3f41;
mem_array[16557] = 16'hf9ca;
mem_array[16556] = 16'hbf8d;
mem_array[16559] = 16'h21d8;
mem_array[16558] = 16'hbfc1;
mem_array[16561] = 16'h91d5;
mem_array[16560] = 16'hbfe2;
mem_array[16563] = 16'h2cf6;
mem_array[16562] = 16'h3e4e;
mem_array[16565] = 16'h8351;
mem_array[16564] = 16'hbf13;
mem_array[16567] = 16'hab69;
mem_array[16566] = 16'hbe90;
mem_array[16569] = 16'h2e0f;
mem_array[16568] = 16'h3ed0;
mem_array[16571] = 16'h1c13;
mem_array[16570] = 16'h3f2f;
mem_array[16573] = 16'h1bc0;
mem_array[16572] = 16'hc043;
mem_array[16575] = 16'h22fc;
mem_array[16574] = 16'h3ddf;
mem_array[16577] = 16'h3983;
mem_array[16576] = 16'hbe29;
mem_array[16579] = 16'h604c;
mem_array[16578] = 16'hbee2;
mem_array[16581] = 16'h1590;
mem_array[16580] = 16'hbda2;
mem_array[16583] = 16'haa71;
mem_array[16582] = 16'h3c7c;
mem_array[16585] = 16'hc095;
mem_array[16584] = 16'hbf91;
mem_array[16587] = 16'h2e87;
mem_array[16586] = 16'hbf87;
mem_array[16589] = 16'ha92a;
mem_array[16588] = 16'h3e62;
mem_array[16591] = 16'h03aa;
mem_array[16590] = 16'hbe93;
mem_array[16593] = 16'he035;
mem_array[16592] = 16'hbefe;
mem_array[16595] = 16'hf75b;
mem_array[16594] = 16'hbf6e;
mem_array[16597] = 16'h3439;
mem_array[16596] = 16'hbe88;
mem_array[16599] = 16'h0cb7;
mem_array[16598] = 16'h3ebf;
mem_array[16601] = 16'h201e;
mem_array[16600] = 16'hbd1e;
mem_array[16603] = 16'h4bc2;
mem_array[16602] = 16'hbd5c;
mem_array[16605] = 16'h5f25;
mem_array[16604] = 16'hbe64;
mem_array[16607] = 16'hf0c8;
mem_array[16606] = 16'hbe9b;
mem_array[16609] = 16'h7a7f;
mem_array[16608] = 16'hbff2;
mem_array[16611] = 16'h2f32;
mem_array[16610] = 16'hbe7a;
mem_array[16613] = 16'h4f91;
mem_array[16612] = 16'h3df0;
mem_array[16615] = 16'h61a0;
mem_array[16614] = 16'h3f95;
mem_array[16617] = 16'h797d;
mem_array[16616] = 16'hbfb9;
mem_array[16619] = 16'ha55b;
mem_array[16618] = 16'hbfbb;
mem_array[16621] = 16'h0a9d;
mem_array[16620] = 16'hbfb6;
mem_array[16623] = 16'h7da8;
mem_array[16622] = 16'h3d9d;
mem_array[16625] = 16'h201f;
mem_array[16624] = 16'hbf04;
mem_array[16627] = 16'h6eac;
mem_array[16626] = 16'hc003;
mem_array[16629] = 16'h32b5;
mem_array[16628] = 16'h3e2c;
mem_array[16631] = 16'h1b33;
mem_array[16630] = 16'h3ed4;
mem_array[16633] = 16'h7e1c;
mem_array[16632] = 16'hbfc3;
mem_array[16635] = 16'hd051;
mem_array[16634] = 16'hbdd0;
mem_array[16637] = 16'h0972;
mem_array[16636] = 16'hbe57;
mem_array[16639] = 16'h089e;
mem_array[16638] = 16'h3c3f;
mem_array[16641] = 16'hedee;
mem_array[16640] = 16'hbd56;
mem_array[16643] = 16'h47a9;
mem_array[16642] = 16'h3cd9;
mem_array[16645] = 16'he4a8;
mem_array[16644] = 16'hbfc6;
mem_array[16647] = 16'hda32;
mem_array[16646] = 16'h3ea4;
mem_array[16649] = 16'ha7e0;
mem_array[16648] = 16'hbf63;
mem_array[16651] = 16'he791;
mem_array[16650] = 16'hbe58;
mem_array[16653] = 16'h1886;
mem_array[16652] = 16'hbe67;
mem_array[16655] = 16'h9349;
mem_array[16654] = 16'h3f7e;
mem_array[16657] = 16'hbaf9;
mem_array[16656] = 16'hbf85;
mem_array[16659] = 16'h8704;
mem_array[16658] = 16'h3efc;
mem_array[16661] = 16'hb520;
mem_array[16660] = 16'hbf59;
mem_array[16663] = 16'hdf09;
mem_array[16662] = 16'h3f36;
mem_array[16665] = 16'h5a38;
mem_array[16664] = 16'hbf36;
mem_array[16667] = 16'h026a;
mem_array[16666] = 16'hbe63;
mem_array[16669] = 16'h1041;
mem_array[16668] = 16'hbf76;
mem_array[16671] = 16'hd034;
mem_array[16670] = 16'hbf80;
mem_array[16673] = 16'h08e1;
mem_array[16672] = 16'h3f8f;
mem_array[16675] = 16'h471a;
mem_array[16674] = 16'h3f3b;
mem_array[16677] = 16'heaa5;
mem_array[16676] = 16'hbf32;
mem_array[16679] = 16'hdfac;
mem_array[16678] = 16'hc00c;
mem_array[16681] = 16'h0d23;
mem_array[16680] = 16'h3fa5;
mem_array[16683] = 16'h24b5;
mem_array[16682] = 16'hbf5f;
mem_array[16685] = 16'h23f8;
mem_array[16684] = 16'hbe22;
mem_array[16687] = 16'h8781;
mem_array[16686] = 16'hbfd4;
mem_array[16689] = 16'h5532;
mem_array[16688] = 16'hbfb4;
mem_array[16691] = 16'h1c3b;
mem_array[16690] = 16'h3f86;
mem_array[16693] = 16'ha363;
mem_array[16692] = 16'h3b62;
mem_array[16695] = 16'h05fd;
mem_array[16694] = 16'h3df9;
mem_array[16697] = 16'ha6f7;
mem_array[16696] = 16'h3ec5;
mem_array[16699] = 16'h488d;
mem_array[16698] = 16'h3e0b;
mem_array[16701] = 16'hf296;
mem_array[16700] = 16'h3d0d;
mem_array[16703] = 16'hd5c7;
mem_array[16702] = 16'h3c89;
mem_array[16705] = 16'h0010;
mem_array[16704] = 16'hbf3b;
mem_array[16707] = 16'h32cc;
mem_array[16706] = 16'hbf4e;
mem_array[16709] = 16'h1aaf;
mem_array[16708] = 16'hbe88;
mem_array[16711] = 16'h38dd;
mem_array[16710] = 16'h3ea7;
mem_array[16713] = 16'h9a89;
mem_array[16712] = 16'hbe8f;
mem_array[16715] = 16'h73aa;
mem_array[16714] = 16'hbf00;
mem_array[16717] = 16'h884d;
mem_array[16716] = 16'hbda8;
mem_array[16719] = 16'h48fc;
mem_array[16718] = 16'h3daa;
mem_array[16721] = 16'hdbfe;
mem_array[16720] = 16'hbf9c;
mem_array[16723] = 16'hbd8d;
mem_array[16722] = 16'hbf11;
mem_array[16725] = 16'h0a0e;
mem_array[16724] = 16'h3e38;
mem_array[16727] = 16'hd729;
mem_array[16726] = 16'hbe81;
mem_array[16729] = 16'h70d6;
mem_array[16728] = 16'hbf84;
mem_array[16731] = 16'hec72;
mem_array[16730] = 16'hbe81;
mem_array[16733] = 16'h1c70;
mem_array[16732] = 16'h3f4e;
mem_array[16735] = 16'he6c6;
mem_array[16734] = 16'h3c0d;
mem_array[16737] = 16'h04b8;
mem_array[16736] = 16'h3f2d;
mem_array[16739] = 16'hdea3;
mem_array[16738] = 16'hbfcc;
mem_array[16741] = 16'hca34;
mem_array[16740] = 16'h3d9d;
mem_array[16743] = 16'h90d9;
mem_array[16742] = 16'hbed1;
mem_array[16745] = 16'h81c6;
mem_array[16744] = 16'hbe74;
mem_array[16747] = 16'hc003;
mem_array[16746] = 16'h3dbf;
mem_array[16749] = 16'ha0ee;
mem_array[16748] = 16'hbe9a;
mem_array[16751] = 16'hf7c0;
mem_array[16750] = 16'h3f75;
mem_array[16753] = 16'h1cfb;
mem_array[16752] = 16'hbd69;
mem_array[16755] = 16'h06ef;
mem_array[16754] = 16'h3de5;
mem_array[16757] = 16'h6027;
mem_array[16756] = 16'h3eb4;
mem_array[16759] = 16'hd99b;
mem_array[16758] = 16'hbe29;
mem_array[16761] = 16'h65de;
mem_array[16760] = 16'h3c92;
mem_array[16763] = 16'hc231;
mem_array[16762] = 16'h3c4f;
mem_array[16765] = 16'hc29e;
mem_array[16764] = 16'hbf71;
mem_array[16767] = 16'hf5d3;
mem_array[16766] = 16'h3d58;
mem_array[16769] = 16'hf4bb;
mem_array[16768] = 16'hbdc2;
mem_array[16771] = 16'hb33c;
mem_array[16770] = 16'h3f1b;
mem_array[16773] = 16'hb5f8;
mem_array[16772] = 16'h3c87;
mem_array[16775] = 16'h34dc;
mem_array[16774] = 16'h3e39;
mem_array[16777] = 16'hbfd5;
mem_array[16776] = 16'hbe3a;
mem_array[16779] = 16'h701e;
mem_array[16778] = 16'hbe73;
mem_array[16781] = 16'hbe27;
mem_array[16780] = 16'hbf30;
mem_array[16783] = 16'h1135;
mem_array[16782] = 16'h3f6b;
mem_array[16785] = 16'hc62b;
mem_array[16784] = 16'h3d76;
mem_array[16787] = 16'h6857;
mem_array[16786] = 16'hbf7e;
mem_array[16789] = 16'h3a04;
mem_array[16788] = 16'hbe12;
mem_array[16791] = 16'h9b1e;
mem_array[16790] = 16'hbeb3;
mem_array[16793] = 16'hb666;
mem_array[16792] = 16'h3f8a;
mem_array[16795] = 16'ha244;
mem_array[16794] = 16'h3f99;
mem_array[16797] = 16'h0cc2;
mem_array[16796] = 16'h3dd8;
mem_array[16799] = 16'h646a;
mem_array[16798] = 16'hbf8c;
mem_array[16801] = 16'h9c72;
mem_array[16800] = 16'hbd3b;
mem_array[16803] = 16'he6a4;
mem_array[16802] = 16'hbd9b;
mem_array[16805] = 16'h4a53;
mem_array[16804] = 16'hbd66;
mem_array[16807] = 16'h3f72;
mem_array[16806] = 16'h3bd4;
mem_array[16809] = 16'h6d70;
mem_array[16808] = 16'h3cf1;
mem_array[16811] = 16'h911a;
mem_array[16810] = 16'hbdd0;
mem_array[16813] = 16'hd7b9;
mem_array[16812] = 16'hbd1d;
mem_array[16815] = 16'ha1c6;
mem_array[16814] = 16'hbd6b;
mem_array[16817] = 16'he9af;
mem_array[16816] = 16'h3d44;
mem_array[16819] = 16'he502;
mem_array[16818] = 16'h3d1a;
mem_array[16821] = 16'h5aed;
mem_array[16820] = 16'hbd92;
mem_array[16823] = 16'h928a;
mem_array[16822] = 16'h3da3;
mem_array[16825] = 16'hcb16;
mem_array[16824] = 16'hbcaa;
mem_array[16827] = 16'h0f56;
mem_array[16826] = 16'h3d25;
mem_array[16829] = 16'he409;
mem_array[16828] = 16'hbdc4;
mem_array[16831] = 16'h3fed;
mem_array[16830] = 16'hbdd3;
mem_array[16833] = 16'h51db;
mem_array[16832] = 16'h3c45;
mem_array[16835] = 16'h40b1;
mem_array[16834] = 16'hbca0;
mem_array[16837] = 16'h987c;
mem_array[16836] = 16'h3db7;
mem_array[16839] = 16'h7ac3;
mem_array[16838] = 16'h3dbf;
mem_array[16841] = 16'h531d;
mem_array[16840] = 16'hbd88;
mem_array[16843] = 16'hd54d;
mem_array[16842] = 16'hb92e;
mem_array[16845] = 16'h3fd2;
mem_array[16844] = 16'hbd68;
mem_array[16847] = 16'h5650;
mem_array[16846] = 16'hbd93;
mem_array[16849] = 16'h80d3;
mem_array[16848] = 16'hbc0b;
mem_array[16851] = 16'hef16;
mem_array[16850] = 16'h3e06;
mem_array[16853] = 16'h1795;
mem_array[16852] = 16'hbe34;
mem_array[16855] = 16'hb070;
mem_array[16854] = 16'h3dec;
mem_array[16857] = 16'h3eec;
mem_array[16856] = 16'h3d04;
mem_array[16859] = 16'h0bf8;
mem_array[16858] = 16'hbd22;
mem_array[16861] = 16'hbbb0;
mem_array[16860] = 16'h3f82;
mem_array[16863] = 16'hc666;
mem_array[16862] = 16'h3f36;
mem_array[16865] = 16'h9ac6;
mem_array[16864] = 16'h3ed1;
mem_array[16867] = 16'h37fd;
mem_array[16866] = 16'hbd1f;
mem_array[16869] = 16'hd418;
mem_array[16868] = 16'hbecf;
mem_array[16871] = 16'hc6b0;
mem_array[16870] = 16'hbcd7;
mem_array[16873] = 16'ha43e;
mem_array[16872] = 16'h3e85;
mem_array[16875] = 16'h94cc;
mem_array[16874] = 16'hbe7d;
mem_array[16877] = 16'hfe33;
mem_array[16876] = 16'hbe31;
mem_array[16879] = 16'h908c;
mem_array[16878] = 16'h3ef6;
mem_array[16881] = 16'he3ac;
mem_array[16880] = 16'hbc33;
mem_array[16883] = 16'hb4d6;
mem_array[16882] = 16'h3d59;
mem_array[16885] = 16'h4c3e;
mem_array[16884] = 16'h3d1b;
mem_array[16887] = 16'hadc0;
mem_array[16886] = 16'h3d55;
mem_array[16889] = 16'heb53;
mem_array[16888] = 16'h3c30;
mem_array[16891] = 16'h9bc6;
mem_array[16890] = 16'hbe3b;
mem_array[16893] = 16'ha6e4;
mem_array[16892] = 16'h3f83;
mem_array[16895] = 16'hbd1a;
mem_array[16894] = 16'h3e98;
mem_array[16897] = 16'h003b;
mem_array[16896] = 16'h3f28;
mem_array[16899] = 16'h41c5;
mem_array[16898] = 16'h3f09;
mem_array[16901] = 16'h7262;
mem_array[16900] = 16'hbeb5;
mem_array[16903] = 16'hb545;
mem_array[16902] = 16'hbe36;
mem_array[16905] = 16'h0eab;
mem_array[16904] = 16'h3dbb;
mem_array[16907] = 16'h9739;
mem_array[16906] = 16'hbf0a;
mem_array[16909] = 16'hc6fd;
mem_array[16908] = 16'hbed7;
mem_array[16911] = 16'hdf73;
mem_array[16910] = 16'h3f03;
mem_array[16913] = 16'h4ad5;
mem_array[16912] = 16'hbf13;
mem_array[16915] = 16'h7a4c;
mem_array[16914] = 16'h3e24;
mem_array[16917] = 16'hed23;
mem_array[16916] = 16'h3e5b;
mem_array[16919] = 16'hc261;
mem_array[16918] = 16'hbf1f;
mem_array[16921] = 16'h3552;
mem_array[16920] = 16'h3db1;
mem_array[16923] = 16'h7b2b;
mem_array[16922] = 16'hbf02;
mem_array[16925] = 16'h94ea;
mem_array[16924] = 16'h3cf6;
mem_array[16927] = 16'h3d2c;
mem_array[16926] = 16'h3e5a;
mem_array[16929] = 16'hcc94;
mem_array[16928] = 16'hbd8d;
mem_array[16931] = 16'he7b8;
mem_array[16930] = 16'hbdbe;
mem_array[16933] = 16'h602d;
mem_array[16932] = 16'h3ecb;
mem_array[16935] = 16'h0be8;
mem_array[16934] = 16'h3e8d;
mem_array[16937] = 16'haa0e;
mem_array[16936] = 16'hbefd;
mem_array[16939] = 16'h15e2;
mem_array[16938] = 16'h3e1d;
mem_array[16941] = 16'h2f7c;
mem_array[16940] = 16'hbce4;
mem_array[16943] = 16'h0fe6;
mem_array[16942] = 16'hbd5b;
mem_array[16945] = 16'hef2f;
mem_array[16944] = 16'hbe66;
mem_array[16947] = 16'he8c5;
mem_array[16946] = 16'h3e02;
mem_array[16949] = 16'hb745;
mem_array[16948] = 16'h3d99;
mem_array[16951] = 16'hc5c3;
mem_array[16950] = 16'hbed8;
mem_array[16953] = 16'hf8c5;
mem_array[16952] = 16'hbef8;
mem_array[16955] = 16'h45f9;
mem_array[16954] = 16'hbe86;
mem_array[16957] = 16'hd09a;
mem_array[16956] = 16'hbe0b;
mem_array[16959] = 16'h0457;
mem_array[16958] = 16'h3eed;
mem_array[16961] = 16'h330e;
mem_array[16960] = 16'hbe9d;
mem_array[16963] = 16'h5901;
mem_array[16962] = 16'h3f04;
mem_array[16965] = 16'h52d3;
mem_array[16964] = 16'h3da9;
mem_array[16967] = 16'h4a82;
mem_array[16966] = 16'h3f8d;
mem_array[16969] = 16'h5228;
mem_array[16968] = 16'hbf1c;
mem_array[16971] = 16'hc95c;
mem_array[16970] = 16'hbe04;
mem_array[16973] = 16'h8b94;
mem_array[16972] = 16'h3df2;
mem_array[16975] = 16'h3d75;
mem_array[16974] = 16'hbb23;
mem_array[16977] = 16'haa4c;
mem_array[16976] = 16'hbdd7;
mem_array[16979] = 16'he9a8;
mem_array[16978] = 16'hbe02;
mem_array[16981] = 16'h93bc;
mem_array[16980] = 16'h3eb2;
mem_array[16983] = 16'hffe4;
mem_array[16982] = 16'hbcba;
mem_array[16985] = 16'hd484;
mem_array[16984] = 16'hbe36;
mem_array[16987] = 16'h25a6;
mem_array[16986] = 16'hbfbe;
mem_array[16989] = 16'hde2d;
mem_array[16988] = 16'h3e34;
mem_array[16991] = 16'hfe3b;
mem_array[16990] = 16'hbed0;
mem_array[16993] = 16'h2c99;
mem_array[16992] = 16'h3f0f;
mem_array[16995] = 16'hd81f;
mem_array[16994] = 16'hbd82;
mem_array[16997] = 16'hf8f5;
mem_array[16996] = 16'hbbe3;
mem_array[16999] = 16'hfc2a;
mem_array[16998] = 16'hbf80;
mem_array[17001] = 16'h1b99;
mem_array[17000] = 16'hbcf3;
mem_array[17003] = 16'h5e0b;
mem_array[17002] = 16'hbd50;
mem_array[17005] = 16'h0fe1;
mem_array[17004] = 16'h3e29;
mem_array[17007] = 16'hab90;
mem_array[17006] = 16'h3e18;
mem_array[17009] = 16'h9b09;
mem_array[17008] = 16'h3e62;
mem_array[17011] = 16'h46b0;
mem_array[17010] = 16'hbda7;
mem_array[17013] = 16'hccd6;
mem_array[17012] = 16'h3e8c;
mem_array[17015] = 16'h398b;
mem_array[17014] = 16'h3f10;
mem_array[17017] = 16'hd48f;
mem_array[17016] = 16'hbda6;
mem_array[17019] = 16'h5f78;
mem_array[17018] = 16'h3e53;
mem_array[17021] = 16'h93bf;
mem_array[17020] = 16'hbeab;
mem_array[17023] = 16'h6cd0;
mem_array[17022] = 16'h3f21;
mem_array[17025] = 16'h0878;
mem_array[17024] = 16'h3e7f;
mem_array[17027] = 16'hdab5;
mem_array[17026] = 16'h3e33;
mem_array[17029] = 16'hc0c4;
mem_array[17028] = 16'h3f4c;
mem_array[17031] = 16'h64b0;
mem_array[17030] = 16'hbf05;
mem_array[17033] = 16'h9879;
mem_array[17032] = 16'h3e76;
mem_array[17035] = 16'he39c;
mem_array[17034] = 16'h3c0b;
mem_array[17037] = 16'h49e8;
mem_array[17036] = 16'hbeb1;
mem_array[17039] = 16'hc1d5;
mem_array[17038] = 16'hbeae;
mem_array[17041] = 16'haf45;
mem_array[17040] = 16'h3f7d;
mem_array[17043] = 16'h62d0;
mem_array[17042] = 16'h3e29;
mem_array[17045] = 16'h3401;
mem_array[17044] = 16'h3da5;
mem_array[17047] = 16'ha9d0;
mem_array[17046] = 16'hbf05;
mem_array[17049] = 16'h3686;
mem_array[17048] = 16'hbf26;
mem_array[17051] = 16'h0fa7;
mem_array[17050] = 16'hbf22;
mem_array[17053] = 16'h07cf;
mem_array[17052] = 16'hbec7;
mem_array[17055] = 16'h4b86;
mem_array[17054] = 16'hbe99;
mem_array[17057] = 16'h36cf;
mem_array[17056] = 16'hbf27;
mem_array[17059] = 16'hd829;
mem_array[17058] = 16'hbe49;
mem_array[17061] = 16'h9790;
mem_array[17060] = 16'hbd52;
mem_array[17063] = 16'h6b0e;
mem_array[17062] = 16'hbd00;
mem_array[17065] = 16'h3331;
mem_array[17064] = 16'h3db8;
mem_array[17067] = 16'h95e2;
mem_array[17066] = 16'h3e88;
mem_array[17069] = 16'h4d58;
mem_array[17068] = 16'hbd10;
mem_array[17071] = 16'h0031;
mem_array[17070] = 16'hbdad;
mem_array[17073] = 16'h742d;
mem_array[17072] = 16'h3f59;
mem_array[17075] = 16'h0919;
mem_array[17074] = 16'h3d09;
mem_array[17077] = 16'h596d;
mem_array[17076] = 16'h3eaa;
mem_array[17079] = 16'h5305;
mem_array[17078] = 16'hbecc;
mem_array[17081] = 16'hb227;
mem_array[17080] = 16'hbef0;
mem_array[17083] = 16'hc7ec;
mem_array[17082] = 16'h3ef0;
mem_array[17085] = 16'hae25;
mem_array[17084] = 16'h3dc8;
mem_array[17087] = 16'hbe5d;
mem_array[17086] = 16'h3dcf;
mem_array[17089] = 16'h38e0;
mem_array[17088] = 16'h3ebd;
mem_array[17091] = 16'h5f89;
mem_array[17090] = 16'h3f27;
mem_array[17093] = 16'hfae6;
mem_array[17092] = 16'h3e82;
mem_array[17095] = 16'hde2b;
mem_array[17094] = 16'hbec5;
mem_array[17097] = 16'h66be;
mem_array[17096] = 16'hbf23;
mem_array[17099] = 16'hec12;
mem_array[17098] = 16'hbed7;
mem_array[17101] = 16'h2046;
mem_array[17100] = 16'h3f1e;
mem_array[17103] = 16'h0941;
mem_array[17102] = 16'h3eb6;
mem_array[17105] = 16'h754e;
mem_array[17104] = 16'h3e54;
mem_array[17107] = 16'hb333;
mem_array[17106] = 16'h3b8b;
mem_array[17109] = 16'h8ffe;
mem_array[17108] = 16'h3e68;
mem_array[17111] = 16'h412f;
mem_array[17110] = 16'hbd50;
mem_array[17113] = 16'h474c;
mem_array[17112] = 16'hbf86;
mem_array[17115] = 16'hfa43;
mem_array[17114] = 16'hbd48;
mem_array[17117] = 16'hd07b;
mem_array[17116] = 16'h3f89;
mem_array[17119] = 16'hd803;
mem_array[17118] = 16'h3e0b;
mem_array[17121] = 16'h0099;
mem_array[17120] = 16'h3dc3;
mem_array[17123] = 16'hd9b5;
mem_array[17122] = 16'hbc50;
mem_array[17125] = 16'he26a;
mem_array[17124] = 16'h3e5a;
mem_array[17127] = 16'h11e2;
mem_array[17126] = 16'h3f0a;
mem_array[17129] = 16'h80e5;
mem_array[17128] = 16'h3e24;
mem_array[17131] = 16'hb928;
mem_array[17130] = 16'hbb89;
mem_array[17133] = 16'h76fc;
mem_array[17132] = 16'h3ee3;
mem_array[17135] = 16'h9a1d;
mem_array[17134] = 16'h3dc7;
mem_array[17137] = 16'hd2a6;
mem_array[17136] = 16'h3c6b;
mem_array[17139] = 16'h6c07;
mem_array[17138] = 16'hbd3a;
mem_array[17141] = 16'h3856;
mem_array[17140] = 16'hbf5b;
mem_array[17143] = 16'h4ec4;
mem_array[17142] = 16'hbd96;
mem_array[17145] = 16'hdc3e;
mem_array[17144] = 16'hbf7b;
mem_array[17147] = 16'h10d8;
mem_array[17146] = 16'hbef6;
mem_array[17149] = 16'hf0e4;
mem_array[17148] = 16'h3ebf;
mem_array[17151] = 16'hed56;
mem_array[17150] = 16'h3ec8;
mem_array[17153] = 16'h6980;
mem_array[17152] = 16'h3d1f;
mem_array[17155] = 16'hddf6;
mem_array[17154] = 16'hbd0f;
mem_array[17157] = 16'h543f;
mem_array[17156] = 16'h3e38;
mem_array[17159] = 16'hce4b;
mem_array[17158] = 16'hbefe;
mem_array[17161] = 16'h20ff;
mem_array[17160] = 16'h3ed1;
mem_array[17163] = 16'hb0d6;
mem_array[17162] = 16'h3d9d;
mem_array[17165] = 16'h4bc1;
mem_array[17164] = 16'h3c9f;
mem_array[17167] = 16'h5a2a;
mem_array[17166] = 16'hbe47;
mem_array[17169] = 16'h3fa6;
mem_array[17168] = 16'h3e16;
mem_array[17171] = 16'h95b2;
mem_array[17170] = 16'hbeeb;
mem_array[17173] = 16'h00f6;
mem_array[17172] = 16'hbf3b;
mem_array[17175] = 16'h4abe;
mem_array[17174] = 16'h3eae;
mem_array[17177] = 16'h9e4c;
mem_array[17176] = 16'h3e58;
mem_array[17179] = 16'h0de3;
mem_array[17178] = 16'hbe4a;
mem_array[17181] = 16'hca83;
mem_array[17180] = 16'hbdfc;
mem_array[17183] = 16'h0059;
mem_array[17182] = 16'h3db0;
mem_array[17185] = 16'h7a73;
mem_array[17184] = 16'h3ed6;
mem_array[17187] = 16'ha1f9;
mem_array[17186] = 16'hbf38;
mem_array[17189] = 16'h5e11;
mem_array[17188] = 16'hbeaf;
mem_array[17191] = 16'h52e2;
mem_array[17190] = 16'h3e45;
mem_array[17193] = 16'h7197;
mem_array[17192] = 16'hbecf;
mem_array[17195] = 16'hcee2;
mem_array[17194] = 16'hbf26;
mem_array[17197] = 16'hfc67;
mem_array[17196] = 16'hbe0d;
mem_array[17199] = 16'hf8f2;
mem_array[17198] = 16'h3da5;
mem_array[17201] = 16'h3f6c;
mem_array[17200] = 16'hbf18;
mem_array[17203] = 16'hfc58;
mem_array[17202] = 16'h3eb1;
mem_array[17205] = 16'h733e;
mem_array[17204] = 16'hbf82;
mem_array[17207] = 16'ha93e;
mem_array[17206] = 16'h3e6a;
mem_array[17209] = 16'h3604;
mem_array[17208] = 16'h3f03;
mem_array[17211] = 16'h7abb;
mem_array[17210] = 16'h3ec5;
mem_array[17213] = 16'h26f6;
mem_array[17212] = 16'h3e5c;
mem_array[17215] = 16'h9690;
mem_array[17214] = 16'hbdb1;
mem_array[17217] = 16'hacb8;
mem_array[17216] = 16'hbeb9;
mem_array[17219] = 16'h6c47;
mem_array[17218] = 16'h3d02;
mem_array[17221] = 16'hca4c;
mem_array[17220] = 16'h3e08;
mem_array[17223] = 16'h9330;
mem_array[17222] = 16'h3ccd;
mem_array[17225] = 16'hd1a5;
mem_array[17224] = 16'hbe65;
mem_array[17227] = 16'h02d9;
mem_array[17226] = 16'hbe9e;
mem_array[17229] = 16'hd39e;
mem_array[17228] = 16'hbe42;
mem_array[17231] = 16'h35e0;
mem_array[17230] = 16'h3e30;
mem_array[17233] = 16'h6fb5;
mem_array[17232] = 16'hbf8b;
mem_array[17235] = 16'hc4b4;
mem_array[17234] = 16'hbeae;
mem_array[17237] = 16'haa98;
mem_array[17236] = 16'h3e5e;
mem_array[17239] = 16'h324e;
mem_array[17238] = 16'h3daf;
mem_array[17241] = 16'h25c3;
mem_array[17240] = 16'hbd28;
mem_array[17243] = 16'hb9f5;
mem_array[17242] = 16'hbdbd;
mem_array[17245] = 16'hd052;
mem_array[17244] = 16'hbd10;
mem_array[17247] = 16'h2eae;
mem_array[17246] = 16'hbf00;
mem_array[17249] = 16'hcd50;
mem_array[17248] = 16'h3e2e;
mem_array[17251] = 16'hb312;
mem_array[17250] = 16'h3e93;
mem_array[17253] = 16'h0d19;
mem_array[17252] = 16'hbe45;
mem_array[17255] = 16'h96ac;
mem_array[17254] = 16'h3b39;
mem_array[17257] = 16'h9ccf;
mem_array[17256] = 16'h3cc1;
mem_array[17259] = 16'h284a;
mem_array[17258] = 16'hbe91;
mem_array[17261] = 16'hb58e;
mem_array[17260] = 16'h3d2c;
mem_array[17263] = 16'hbdac;
mem_array[17262] = 16'h3e84;
mem_array[17265] = 16'h551f;
mem_array[17264] = 16'hbe02;
mem_array[17267] = 16'hdaae;
mem_array[17266] = 16'h3e8a;
mem_array[17269] = 16'h0bf0;
mem_array[17268] = 16'h3ebe;
mem_array[17271] = 16'h14ec;
mem_array[17270] = 16'h3ab8;
mem_array[17273] = 16'h2dfe;
mem_array[17272] = 16'h3d5e;
mem_array[17275] = 16'h9ebd;
mem_array[17274] = 16'hbe85;
mem_array[17277] = 16'hd602;
mem_array[17276] = 16'hbf2d;
mem_array[17279] = 16'hdf21;
mem_array[17278] = 16'hbed3;
mem_array[17281] = 16'h0bf0;
mem_array[17280] = 16'h3d6b;
mem_array[17283] = 16'hef23;
mem_array[17282] = 16'hbd86;
mem_array[17285] = 16'h25e5;
mem_array[17284] = 16'h3e1a;
mem_array[17287] = 16'h8f1c;
mem_array[17286] = 16'hbe9a;
mem_array[17289] = 16'h2f81;
mem_array[17288] = 16'hbe0e;
mem_array[17291] = 16'had8c;
mem_array[17290] = 16'hbc99;
mem_array[17293] = 16'hb9e9;
mem_array[17292] = 16'hbffc;
mem_array[17295] = 16'hab59;
mem_array[17294] = 16'hbedd;
mem_array[17297] = 16'h128e;
mem_array[17296] = 16'h3df5;
mem_array[17299] = 16'he935;
mem_array[17298] = 16'hbe8e;
mem_array[17301] = 16'h5bc0;
mem_array[17300] = 16'hbd79;
mem_array[17303] = 16'h46f3;
mem_array[17302] = 16'h3d29;
mem_array[17305] = 16'h8bea;
mem_array[17304] = 16'hbe9f;
mem_array[17307] = 16'h8312;
mem_array[17306] = 16'h3e18;
mem_array[17309] = 16'hd36e;
mem_array[17308] = 16'h3e64;
mem_array[17311] = 16'h0329;
mem_array[17310] = 16'h3c56;
mem_array[17313] = 16'h925e;
mem_array[17312] = 16'hbe71;
mem_array[17315] = 16'h1b85;
mem_array[17314] = 16'h3d36;
mem_array[17317] = 16'h6306;
mem_array[17316] = 16'h3d9b;
mem_array[17319] = 16'ha294;
mem_array[17318] = 16'hbd19;
mem_array[17321] = 16'h0e83;
mem_array[17320] = 16'h3e3b;
mem_array[17323] = 16'hcbf8;
mem_array[17322] = 16'h3e3f;
mem_array[17325] = 16'h8880;
mem_array[17324] = 16'hbf0e;
mem_array[17327] = 16'hea84;
mem_array[17326] = 16'hbd1c;
mem_array[17329] = 16'h84b6;
mem_array[17328] = 16'h3f59;
mem_array[17331] = 16'hd533;
mem_array[17330] = 16'hb9f4;
mem_array[17333] = 16'h8f40;
mem_array[17332] = 16'h3d8f;
mem_array[17335] = 16'heaf3;
mem_array[17334] = 16'h3e13;
mem_array[17337] = 16'haae7;
mem_array[17336] = 16'hbf61;
mem_array[17339] = 16'h9b0f;
mem_array[17338] = 16'hbeb8;
mem_array[17341] = 16'h3c24;
mem_array[17340] = 16'hbe0e;
mem_array[17343] = 16'h251d;
mem_array[17342] = 16'hbc57;
mem_array[17345] = 16'hdf54;
mem_array[17344] = 16'h3c30;
mem_array[17347] = 16'ha977;
mem_array[17346] = 16'hbdd7;
mem_array[17349] = 16'h0899;
mem_array[17348] = 16'hbe02;
mem_array[17351] = 16'ha349;
mem_array[17350] = 16'h3cfd;
mem_array[17353] = 16'hc497;
mem_array[17352] = 16'hbff1;
mem_array[17355] = 16'ha944;
mem_array[17354] = 16'h3e8c;
mem_array[17357] = 16'hc011;
mem_array[17356] = 16'h3e99;
mem_array[17359] = 16'hf371;
mem_array[17358] = 16'hbeba;
mem_array[17361] = 16'hede9;
mem_array[17360] = 16'hbe00;
mem_array[17363] = 16'hc44f;
mem_array[17362] = 16'hbd9d;
mem_array[17365] = 16'he4b7;
mem_array[17364] = 16'hbe67;
mem_array[17367] = 16'h397a;
mem_array[17366] = 16'h3e64;
mem_array[17369] = 16'ha461;
mem_array[17368] = 16'hbdbe;
mem_array[17371] = 16'h14d5;
mem_array[17370] = 16'hbde2;
mem_array[17373] = 16'hf5b2;
mem_array[17372] = 16'h3d35;
mem_array[17375] = 16'h2ea6;
mem_array[17374] = 16'hbd1c;
mem_array[17377] = 16'hf41d;
mem_array[17376] = 16'h3e58;
mem_array[17379] = 16'hf01e;
mem_array[17378] = 16'hbe04;
mem_array[17381] = 16'hc7ea;
mem_array[17380] = 16'hbe42;
mem_array[17383] = 16'hc4b0;
mem_array[17382] = 16'h3e2e;
mem_array[17385] = 16'hf11c;
mem_array[17384] = 16'hbe68;
mem_array[17387] = 16'hc794;
mem_array[17386] = 16'h3c10;
mem_array[17389] = 16'hf0b8;
mem_array[17388] = 16'h3ef2;
mem_array[17391] = 16'h0bee;
mem_array[17390] = 16'h3eb3;
mem_array[17393] = 16'hbece;
mem_array[17392] = 16'h3e20;
mem_array[17395] = 16'h745d;
mem_array[17394] = 16'hbda0;
mem_array[17397] = 16'h8775;
mem_array[17396] = 16'hbf2d;
mem_array[17399] = 16'h83a7;
mem_array[17398] = 16'hbefe;
mem_array[17401] = 16'h42f8;
mem_array[17400] = 16'hbea3;
mem_array[17403] = 16'h1b6c;
mem_array[17402] = 16'h3ca8;
mem_array[17405] = 16'h5c0d;
mem_array[17404] = 16'hbd2a;
mem_array[17407] = 16'hfc65;
mem_array[17406] = 16'hbeb8;
mem_array[17409] = 16'h5f8e;
mem_array[17408] = 16'h3c05;
mem_array[17411] = 16'h9e9b;
mem_array[17410] = 16'h3cb7;
mem_array[17413] = 16'h232c;
mem_array[17412] = 16'hbf8a;
mem_array[17415] = 16'h7ac4;
mem_array[17414] = 16'h3eb7;
mem_array[17417] = 16'hb948;
mem_array[17416] = 16'h3e6b;
mem_array[17419] = 16'hc106;
mem_array[17418] = 16'hbc05;
mem_array[17421] = 16'h3fa8;
mem_array[17420] = 16'hbc5c;
mem_array[17423] = 16'h3976;
mem_array[17422] = 16'h3b99;
mem_array[17425] = 16'h777d;
mem_array[17424] = 16'hbebe;
mem_array[17427] = 16'he1b3;
mem_array[17426] = 16'hbe9b;
mem_array[17429] = 16'hebcf;
mem_array[17428] = 16'hbe0f;
mem_array[17431] = 16'h776e;
mem_array[17430] = 16'h3df9;
mem_array[17433] = 16'hb11b;
mem_array[17432] = 16'hbf16;
mem_array[17435] = 16'h2e6e;
mem_array[17434] = 16'h3c03;
mem_array[17437] = 16'h222d;
mem_array[17436] = 16'hbe12;
mem_array[17439] = 16'hf3a5;
mem_array[17438] = 16'hbd9a;
mem_array[17441] = 16'h1e6d;
mem_array[17440] = 16'h3d5e;
mem_array[17443] = 16'hc18d;
mem_array[17442] = 16'h3da1;
mem_array[17445] = 16'he03c;
mem_array[17444] = 16'hbe84;
mem_array[17447] = 16'h340a;
mem_array[17446] = 16'hbd03;
mem_array[17449] = 16'hfcb0;
mem_array[17448] = 16'h3edb;
mem_array[17451] = 16'hb7b4;
mem_array[17450] = 16'h3e31;
mem_array[17453] = 16'h80cb;
mem_array[17452] = 16'h3cb1;
mem_array[17455] = 16'h8d43;
mem_array[17454] = 16'h3e4e;
mem_array[17457] = 16'h9cd1;
mem_array[17456] = 16'hbead;
mem_array[17459] = 16'h5d83;
mem_array[17458] = 16'hbf28;
mem_array[17461] = 16'h6742;
mem_array[17460] = 16'hbf0c;
mem_array[17463] = 16'h4483;
mem_array[17462] = 16'h3f3d;
mem_array[17465] = 16'h6349;
mem_array[17464] = 16'hbe07;
mem_array[17467] = 16'h42f2;
mem_array[17466] = 16'hbe8c;
mem_array[17469] = 16'hea42;
mem_array[17468] = 16'hbe28;
mem_array[17471] = 16'h3971;
mem_array[17470] = 16'h3df7;
mem_array[17473] = 16'h9f8c;
mem_array[17472] = 16'hbf28;
mem_array[17475] = 16'hfa3d;
mem_array[17474] = 16'h3d59;
mem_array[17477] = 16'h39ce;
mem_array[17476] = 16'h3ea0;
mem_array[17479] = 16'hd9d4;
mem_array[17478] = 16'hbe5c;
mem_array[17481] = 16'h2922;
mem_array[17480] = 16'hbb69;
mem_array[17483] = 16'h205b;
mem_array[17482] = 16'h3d05;
mem_array[17485] = 16'h7225;
mem_array[17484] = 16'hbeb4;
mem_array[17487] = 16'hc1f4;
mem_array[17486] = 16'hbedb;
mem_array[17489] = 16'hd5bc;
mem_array[17488] = 16'h3e0f;
mem_array[17491] = 16'h2a09;
mem_array[17490] = 16'hbd53;
mem_array[17493] = 16'h0902;
mem_array[17492] = 16'hbf7e;
mem_array[17495] = 16'heb5c;
mem_array[17494] = 16'hbb1a;
mem_array[17497] = 16'h1905;
mem_array[17496] = 16'h3dbc;
mem_array[17499] = 16'h4f35;
mem_array[17498] = 16'hbe12;
mem_array[17501] = 16'h984e;
mem_array[17500] = 16'hbe15;
mem_array[17503] = 16'h4e87;
mem_array[17502] = 16'h3d52;
mem_array[17505] = 16'ha41e;
mem_array[17504] = 16'hbda8;
mem_array[17507] = 16'h1649;
mem_array[17506] = 16'hbdf5;
mem_array[17509] = 16'h36d4;
mem_array[17508] = 16'hbe5d;
mem_array[17511] = 16'h2d9b;
mem_array[17510] = 16'h3e60;
mem_array[17513] = 16'h962b;
mem_array[17512] = 16'hbe3c;
mem_array[17515] = 16'hc65a;
mem_array[17514] = 16'h3e89;
mem_array[17517] = 16'h9851;
mem_array[17516] = 16'hbeb1;
mem_array[17519] = 16'ha359;
mem_array[17518] = 16'hbe20;
mem_array[17521] = 16'h1c64;
mem_array[17520] = 16'hbecf;
mem_array[17523] = 16'hd253;
mem_array[17522] = 16'h3e39;
mem_array[17525] = 16'hae38;
mem_array[17524] = 16'hbd67;
mem_array[17527] = 16'h8c21;
mem_array[17526] = 16'h3db6;
mem_array[17529] = 16'h90cb;
mem_array[17528] = 16'hbe60;
mem_array[17531] = 16'h80f3;
mem_array[17530] = 16'hbc21;
mem_array[17533] = 16'h87f4;
mem_array[17532] = 16'hbeb4;
mem_array[17535] = 16'h041c;
mem_array[17534] = 16'hbdc3;
mem_array[17537] = 16'h3828;
mem_array[17536] = 16'h3e14;
mem_array[17539] = 16'hcf06;
mem_array[17538] = 16'hbee0;
mem_array[17541] = 16'h6e73;
mem_array[17540] = 16'hbd9a;
mem_array[17543] = 16'hb1df;
mem_array[17542] = 16'h3c4e;
mem_array[17545] = 16'h07e6;
mem_array[17544] = 16'hbf18;
mem_array[17547] = 16'h7374;
mem_array[17546] = 16'hbe09;
mem_array[17549] = 16'h12e7;
mem_array[17548] = 16'h3ec8;
mem_array[17551] = 16'had36;
mem_array[17550] = 16'h3e56;
mem_array[17553] = 16'hc5c3;
mem_array[17552] = 16'hbe2a;
mem_array[17555] = 16'hc7c7;
mem_array[17554] = 16'h3ecc;
mem_array[17557] = 16'ha23f;
mem_array[17556] = 16'h3d66;
mem_array[17559] = 16'hcab9;
mem_array[17558] = 16'h3e2f;
mem_array[17561] = 16'h7a7c;
mem_array[17560] = 16'hbd37;
mem_array[17563] = 16'hb7ff;
mem_array[17562] = 16'h3e7c;
mem_array[17565] = 16'h1458;
mem_array[17564] = 16'hbe81;
mem_array[17567] = 16'hbf9c;
mem_array[17566] = 16'h3e7d;
mem_array[17569] = 16'hc2eb;
mem_array[17568] = 16'hbf0f;
mem_array[17571] = 16'he20d;
mem_array[17570] = 16'h3d5a;
mem_array[17573] = 16'h6f7c;
mem_array[17572] = 16'hbd3a;
mem_array[17575] = 16'h5302;
mem_array[17574] = 16'h3d87;
mem_array[17577] = 16'h1293;
mem_array[17576] = 16'hbe87;
mem_array[17579] = 16'h49d4;
mem_array[17578] = 16'hbc8f;
mem_array[17581] = 16'hc61a;
mem_array[17580] = 16'hbf3d;
mem_array[17583] = 16'h6b6f;
mem_array[17582] = 16'h3dca;
mem_array[17585] = 16'h6d05;
mem_array[17584] = 16'hbec8;
mem_array[17587] = 16'h37ed;
mem_array[17586] = 16'hbe8e;
mem_array[17589] = 16'h4523;
mem_array[17588] = 16'hbd91;
mem_array[17591] = 16'hc41c;
mem_array[17590] = 16'h3e99;
mem_array[17593] = 16'hd415;
mem_array[17592] = 16'h3ee7;
mem_array[17595] = 16'ha98f;
mem_array[17594] = 16'h3e86;
mem_array[17597] = 16'hff5c;
mem_array[17596] = 16'hbe1d;
mem_array[17599] = 16'h517b;
mem_array[17598] = 16'h3f3e;
mem_array[17601] = 16'h56f1;
mem_array[17600] = 16'hbcf7;
mem_array[17603] = 16'h7aa7;
mem_array[17602] = 16'hbc0a;
mem_array[17605] = 16'h37fd;
mem_array[17604] = 16'hbe84;
mem_array[17607] = 16'he1e4;
mem_array[17606] = 16'hbf49;
mem_array[17609] = 16'h06c2;
mem_array[17608] = 16'h3ec5;
mem_array[17611] = 16'hf532;
mem_array[17610] = 16'hbe20;
mem_array[17613] = 16'hfa1c;
mem_array[17612] = 16'hbe88;
mem_array[17615] = 16'h303b;
mem_array[17614] = 16'hbf26;
mem_array[17617] = 16'hd2c3;
mem_array[17616] = 16'hbdc5;
mem_array[17619] = 16'haf0c;
mem_array[17618] = 16'h3dc1;
mem_array[17621] = 16'hf76b;
mem_array[17620] = 16'hbe10;
mem_array[17623] = 16'hb5bf;
mem_array[17622] = 16'h3e47;
mem_array[17625] = 16'h29d9;
mem_array[17624] = 16'hbe28;
mem_array[17627] = 16'h9f6e;
mem_array[17626] = 16'h3daf;
mem_array[17629] = 16'h1146;
mem_array[17628] = 16'hbfa3;
mem_array[17631] = 16'h4cda;
mem_array[17630] = 16'h3cda;
mem_array[17633] = 16'h41ea;
mem_array[17632] = 16'hbe9e;
mem_array[17635] = 16'hb2a6;
mem_array[17634] = 16'h3ea2;
mem_array[17637] = 16'h22ec;
mem_array[17636] = 16'hbf17;
mem_array[17639] = 16'hc23f;
mem_array[17638] = 16'hbdb0;
mem_array[17641] = 16'hf331;
mem_array[17640] = 16'hbe1c;
mem_array[17643] = 16'hdbe3;
mem_array[17642] = 16'hbe1d;
mem_array[17645] = 16'h00ad;
mem_array[17644] = 16'hbf5a;
mem_array[17647] = 16'hb47c;
mem_array[17646] = 16'h3ec8;
mem_array[17649] = 16'h32b2;
mem_array[17648] = 16'hbf28;
mem_array[17651] = 16'h631e;
mem_array[17650] = 16'h3bb6;
mem_array[17653] = 16'h97a0;
mem_array[17652] = 16'h3f00;
mem_array[17655] = 16'hdfa6;
mem_array[17654] = 16'h3db6;
mem_array[17657] = 16'hdb3f;
mem_array[17656] = 16'h3e49;
mem_array[17659] = 16'h88ad;
mem_array[17658] = 16'h3f1b;
mem_array[17661] = 16'h7662;
mem_array[17660] = 16'hbcfa;
mem_array[17663] = 16'hd644;
mem_array[17662] = 16'h3d3b;
mem_array[17665] = 16'h56bd;
mem_array[17664] = 16'hbd69;
mem_array[17667] = 16'h169c;
mem_array[17666] = 16'hbeea;
mem_array[17669] = 16'hc663;
mem_array[17668] = 16'hbea6;
mem_array[17671] = 16'ha353;
mem_array[17670] = 16'h3e30;
mem_array[17673] = 16'hf1ae;
mem_array[17672] = 16'h3ea4;
mem_array[17675] = 16'hc1f8;
mem_array[17674] = 16'hbff7;
mem_array[17677] = 16'h8c10;
mem_array[17676] = 16'hbd46;
mem_array[17679] = 16'h65b3;
mem_array[17678] = 16'hbf23;
mem_array[17681] = 16'h0d27;
mem_array[17680] = 16'hbe23;
mem_array[17683] = 16'h7456;
mem_array[17682] = 16'h3e9b;
mem_array[17685] = 16'h6771;
mem_array[17684] = 16'hbea8;
mem_array[17687] = 16'h47e1;
mem_array[17686] = 16'h3e31;
mem_array[17689] = 16'h9781;
mem_array[17688] = 16'hbf62;
mem_array[17691] = 16'h064e;
mem_array[17690] = 16'hbefb;
mem_array[17693] = 16'h496a;
mem_array[17692] = 16'hbeaf;
mem_array[17695] = 16'h56af;
mem_array[17694] = 16'h3d7a;
mem_array[17697] = 16'h9447;
mem_array[17696] = 16'h3cfe;
mem_array[17699] = 16'hea48;
mem_array[17698] = 16'hbdfb;
mem_array[17701] = 16'h0ffe;
mem_array[17700] = 16'h3ec1;
mem_array[17703] = 16'had84;
mem_array[17702] = 16'hbdd4;
mem_array[17705] = 16'h2fb2;
mem_array[17704] = 16'hbed1;
mem_array[17707] = 16'h44b4;
mem_array[17706] = 16'h3e88;
mem_array[17709] = 16'hf4f1;
mem_array[17708] = 16'hbea0;
mem_array[17711] = 16'hd13d;
mem_array[17710] = 16'hbeaa;
mem_array[17713] = 16'h7ead;
mem_array[17712] = 16'h3e5c;
mem_array[17715] = 16'h7eaa;
mem_array[17714] = 16'h3b02;
mem_array[17717] = 16'he122;
mem_array[17716] = 16'h3e97;
mem_array[17719] = 16'ha471;
mem_array[17718] = 16'h3ef1;
mem_array[17721] = 16'he5be;
mem_array[17720] = 16'hbe13;
mem_array[17723] = 16'h6a07;
mem_array[17722] = 16'hbdcc;
mem_array[17725] = 16'hc948;
mem_array[17724] = 16'h3d32;
mem_array[17727] = 16'h2ff9;
mem_array[17726] = 16'hbf2c;
mem_array[17729] = 16'hdb9e;
mem_array[17728] = 16'hbf24;
mem_array[17731] = 16'h4299;
mem_array[17730] = 16'h3dd6;
mem_array[17733] = 16'hcaa7;
mem_array[17732] = 16'h3d8b;
mem_array[17735] = 16'hde14;
mem_array[17734] = 16'hbe3a;
mem_array[17737] = 16'he73b;
mem_array[17736] = 16'h3d8e;
mem_array[17739] = 16'h2793;
mem_array[17738] = 16'hbf5a;
mem_array[17741] = 16'hb355;
mem_array[17740] = 16'h3e8e;
mem_array[17743] = 16'he46d;
mem_array[17742] = 16'h3c9c;
mem_array[17745] = 16'hdab6;
mem_array[17744] = 16'hbe97;
mem_array[17747] = 16'h3874;
mem_array[17746] = 16'h3d23;
mem_array[17749] = 16'h2e80;
mem_array[17748] = 16'hbd97;
mem_array[17751] = 16'h307f;
mem_array[17750] = 16'h3dc2;
mem_array[17753] = 16'h8123;
mem_array[17752] = 16'hbef5;
mem_array[17755] = 16'h3168;
mem_array[17754] = 16'h3e19;
mem_array[17757] = 16'h15b3;
mem_array[17756] = 16'h3e89;
mem_array[17759] = 16'h04bb;
mem_array[17758] = 16'h3e0d;
mem_array[17761] = 16'hb11f;
mem_array[17760] = 16'h3f17;
mem_array[17763] = 16'hb1f9;
mem_array[17762] = 16'hbe09;
mem_array[17765] = 16'h0bc4;
mem_array[17764] = 16'hbbab;
mem_array[17767] = 16'h6595;
mem_array[17766] = 16'hbd5b;
mem_array[17769] = 16'hf51b;
mem_array[17768] = 16'hbe46;
mem_array[17771] = 16'h3d5b;
mem_array[17770] = 16'hbf6e;
mem_array[17773] = 16'ha632;
mem_array[17772] = 16'h3e10;
mem_array[17775] = 16'h148f;
mem_array[17774] = 16'h3d88;
mem_array[17777] = 16'h2943;
mem_array[17776] = 16'h3eb6;
mem_array[17779] = 16'hd93b;
mem_array[17778] = 16'h3d2e;
mem_array[17781] = 16'h8cf8;
mem_array[17780] = 16'hbd2b;
mem_array[17783] = 16'h1057;
mem_array[17782] = 16'hbda3;
mem_array[17785] = 16'hd4e0;
mem_array[17784] = 16'h3e08;
mem_array[17787] = 16'h96ce;
mem_array[17786] = 16'hbdce;
mem_array[17789] = 16'hd56b;
mem_array[17788] = 16'hbef5;
mem_array[17791] = 16'h7db7;
mem_array[17790] = 16'h3e9d;
mem_array[17793] = 16'h18f8;
mem_array[17792] = 16'h3e76;
mem_array[17795] = 16'h92f7;
mem_array[17794] = 16'h3ded;
mem_array[17797] = 16'h8e67;
mem_array[17796] = 16'h3ea0;
mem_array[17799] = 16'h3e79;
mem_array[17798] = 16'hbdd4;
mem_array[17801] = 16'hd8a6;
mem_array[17800] = 16'hbe1f;
mem_array[17803] = 16'hce53;
mem_array[17802] = 16'hbc00;
mem_array[17805] = 16'hcc48;
mem_array[17804] = 16'hbf92;
mem_array[17807] = 16'h9a98;
mem_array[17806] = 16'hbd02;
mem_array[17809] = 16'h2d20;
mem_array[17808] = 16'h3b9d;
mem_array[17811] = 16'h8e44;
mem_array[17810] = 16'h3e8a;
mem_array[17813] = 16'he7af;
mem_array[17812] = 16'hbef0;
mem_array[17815] = 16'h0ae0;
mem_array[17814] = 16'h3e4d;
mem_array[17817] = 16'h7f78;
mem_array[17816] = 16'h3d8d;
mem_array[17819] = 16'h3880;
mem_array[17818] = 16'h3db6;
mem_array[17821] = 16'he682;
mem_array[17820] = 16'h3ec0;
mem_array[17823] = 16'h4e25;
mem_array[17822] = 16'hbe09;
mem_array[17825] = 16'hf4c3;
mem_array[17824] = 16'h3d54;
mem_array[17827] = 16'hcf91;
mem_array[17826] = 16'h3e24;
mem_array[17829] = 16'hcebd;
mem_array[17828] = 16'h3e92;
mem_array[17831] = 16'hcfae;
mem_array[17830] = 16'hbf9d;
mem_array[17833] = 16'h84d9;
mem_array[17832] = 16'hbba2;
mem_array[17835] = 16'h1225;
mem_array[17834] = 16'hbdf9;
mem_array[17837] = 16'hbe18;
mem_array[17836] = 16'h3e1f;
mem_array[17839] = 16'hf9c3;
mem_array[17838] = 16'hbdd4;
mem_array[17841] = 16'h6a95;
mem_array[17840] = 16'h3c59;
mem_array[17843] = 16'h302b;
mem_array[17842] = 16'h3cad;
mem_array[17845] = 16'h9bef;
mem_array[17844] = 16'h3eea;
mem_array[17847] = 16'h4173;
mem_array[17846] = 16'hbdc7;
mem_array[17849] = 16'h11a0;
mem_array[17848] = 16'hbd2a;
mem_array[17851] = 16'hcc55;
mem_array[17850] = 16'h3ee4;
mem_array[17853] = 16'h0eec;
mem_array[17852] = 16'h3e90;
mem_array[17855] = 16'h2ef7;
mem_array[17854] = 16'h3e7c;
mem_array[17857] = 16'hd36f;
mem_array[17856] = 16'h3d7a;
mem_array[17859] = 16'h98aa;
mem_array[17858] = 16'h3ef3;
mem_array[17861] = 16'h5971;
mem_array[17860] = 16'h3bb7;
mem_array[17863] = 16'hdb39;
mem_array[17862] = 16'h3c84;
mem_array[17865] = 16'h4de6;
mem_array[17864] = 16'hbf9b;
mem_array[17867] = 16'h89e4;
mem_array[17866] = 16'h3e24;
mem_array[17869] = 16'hdf39;
mem_array[17868] = 16'hbce0;
mem_array[17871] = 16'hc20e;
mem_array[17870] = 16'h3e94;
mem_array[17873] = 16'h96b5;
mem_array[17872] = 16'hbf05;
mem_array[17875] = 16'h83ef;
mem_array[17874] = 16'h3e80;
mem_array[17877] = 16'h0741;
mem_array[17876] = 16'h3d8a;
mem_array[17879] = 16'h042c;
mem_array[17878] = 16'hbd68;
mem_array[17881] = 16'hfd73;
mem_array[17880] = 16'h3e27;
mem_array[17883] = 16'h8f39;
mem_array[17882] = 16'h3e0f;
mem_array[17885] = 16'h9280;
mem_array[17884] = 16'h3e05;
mem_array[17887] = 16'hef90;
mem_array[17886] = 16'h3e89;
mem_array[17889] = 16'h7cea;
mem_array[17888] = 16'h3dae;
mem_array[17891] = 16'h0efd;
mem_array[17890] = 16'hc00c;
mem_array[17893] = 16'hb3da;
mem_array[17892] = 16'h3d41;
mem_array[17895] = 16'hd238;
mem_array[17894] = 16'hbe8a;
mem_array[17897] = 16'h8f92;
mem_array[17896] = 16'hbca3;
mem_array[17899] = 16'h230b;
mem_array[17898] = 16'hbea2;
mem_array[17901] = 16'h8355;
mem_array[17900] = 16'h3c09;
mem_array[17903] = 16'hbdc9;
mem_array[17902] = 16'hbca5;
mem_array[17905] = 16'h29cb;
mem_array[17904] = 16'hbd14;
mem_array[17907] = 16'h79b8;
mem_array[17906] = 16'hbb9b;
mem_array[17909] = 16'h9dac;
mem_array[17908] = 16'h3e03;
mem_array[17911] = 16'h4022;
mem_array[17910] = 16'h3ed8;
mem_array[17913] = 16'he919;
mem_array[17912] = 16'h3dbe;
mem_array[17915] = 16'hd7bc;
mem_array[17914] = 16'hbc1b;
mem_array[17917] = 16'h82a7;
mem_array[17916] = 16'h3ce2;
mem_array[17919] = 16'h20bc;
mem_array[17918] = 16'h3e69;
mem_array[17921] = 16'hdd54;
mem_array[17920] = 16'h3d77;
mem_array[17923] = 16'h77fd;
mem_array[17922] = 16'hbda9;
mem_array[17925] = 16'hd1f6;
mem_array[17924] = 16'hbfc5;
mem_array[17927] = 16'ha44f;
mem_array[17926] = 16'h3d19;
mem_array[17929] = 16'he3ef;
mem_array[17928] = 16'h3e15;
mem_array[17931] = 16'h4e9e;
mem_array[17930] = 16'h3def;
mem_array[17933] = 16'heda0;
mem_array[17932] = 16'hbe7b;
mem_array[17935] = 16'h76cd;
mem_array[17934] = 16'h3e8f;
mem_array[17937] = 16'h3f6a;
mem_array[17936] = 16'h3e2b;
mem_array[17939] = 16'h0526;
mem_array[17938] = 16'hbe89;
mem_array[17941] = 16'hd597;
mem_array[17940] = 16'hbddb;
mem_array[17943] = 16'h9a4b;
mem_array[17942] = 16'h3e53;
mem_array[17945] = 16'hd447;
mem_array[17944] = 16'hbe35;
mem_array[17947] = 16'h713e;
mem_array[17946] = 16'h3e15;
mem_array[17949] = 16'hb4e7;
mem_array[17948] = 16'h3e93;
mem_array[17951] = 16'h8d1b;
mem_array[17950] = 16'hbfd0;
mem_array[17953] = 16'h2959;
mem_array[17952] = 16'h3e29;
mem_array[17955] = 16'h2bd0;
mem_array[17954] = 16'h3dfc;
mem_array[17957] = 16'hfd81;
mem_array[17956] = 16'hbe52;
mem_array[17959] = 16'hbd13;
mem_array[17958] = 16'hbf92;
mem_array[17961] = 16'h0546;
mem_array[17960] = 16'hbe2e;
mem_array[17963] = 16'h07a7;
mem_array[17962] = 16'h3c92;
mem_array[17965] = 16'h618c;
mem_array[17964] = 16'hbd7b;
mem_array[17967] = 16'hcebe;
mem_array[17966] = 16'hbdc7;
mem_array[17969] = 16'hcd73;
mem_array[17968] = 16'h3e02;
mem_array[17971] = 16'h975a;
mem_array[17970] = 16'h3ef1;
mem_array[17973] = 16'hafe2;
mem_array[17972] = 16'hbd9f;
mem_array[17975] = 16'h990d;
mem_array[17974] = 16'h3e28;
mem_array[17977] = 16'h803a;
mem_array[17976] = 16'hbcec;
mem_array[17979] = 16'h3c6e;
mem_array[17978] = 16'h3e2a;
mem_array[17981] = 16'h1bbf;
mem_array[17980] = 16'hbd0d;
mem_array[17983] = 16'hdb40;
mem_array[17982] = 16'hbd89;
mem_array[17985] = 16'ha48e;
mem_array[17984] = 16'hbfb7;
mem_array[17987] = 16'h6000;
mem_array[17986] = 16'hbc60;
mem_array[17989] = 16'h58f1;
mem_array[17988] = 16'h3cc2;
mem_array[17991] = 16'h0b61;
mem_array[17990] = 16'h3e64;
mem_array[17993] = 16'h20d2;
mem_array[17992] = 16'hbe95;
mem_array[17995] = 16'h6dd3;
mem_array[17994] = 16'h3edb;
mem_array[17997] = 16'hb5fb;
mem_array[17996] = 16'h3e7d;
mem_array[17999] = 16'hbd41;
mem_array[17998] = 16'hbebc;
mem_array[18001] = 16'he3d8;
mem_array[18000] = 16'hbee1;
mem_array[18003] = 16'hf581;
mem_array[18002] = 16'h3dab;
mem_array[18005] = 16'h0968;
mem_array[18004] = 16'hbd9c;
mem_array[18007] = 16'h9e1a;
mem_array[18006] = 16'h3e54;
mem_array[18009] = 16'hfd84;
mem_array[18008] = 16'hbc91;
mem_array[18011] = 16'h08d5;
mem_array[18010] = 16'hbf14;
mem_array[18013] = 16'h08a9;
mem_array[18012] = 16'hbe23;
mem_array[18015] = 16'h56df;
mem_array[18014] = 16'hbd94;
mem_array[18017] = 16'h85bb;
mem_array[18016] = 16'hbed9;
mem_array[18019] = 16'h0aec;
mem_array[18018] = 16'hbf7d;
mem_array[18021] = 16'h213b;
mem_array[18020] = 16'hbd97;
mem_array[18023] = 16'h2d7e;
mem_array[18022] = 16'h3b8f;
mem_array[18025] = 16'h9a3f;
mem_array[18024] = 16'h3d90;
mem_array[18027] = 16'h331d;
mem_array[18026] = 16'hbe83;
mem_array[18029] = 16'hecd0;
mem_array[18028] = 16'h3e87;
mem_array[18031] = 16'h5ecc;
mem_array[18030] = 16'h3e5c;
mem_array[18033] = 16'h0f43;
mem_array[18032] = 16'hbe58;
mem_array[18035] = 16'h9fdc;
mem_array[18034] = 16'hbe25;
mem_array[18037] = 16'h518f;
mem_array[18036] = 16'hbd50;
mem_array[18039] = 16'h3139;
mem_array[18038] = 16'h3e5a;
mem_array[18041] = 16'h7b45;
mem_array[18040] = 16'h3e03;
mem_array[18043] = 16'h091a;
mem_array[18042] = 16'hbe5b;
mem_array[18045] = 16'h20a6;
mem_array[18044] = 16'hbe52;
mem_array[18047] = 16'h5032;
mem_array[18046] = 16'h3c77;
mem_array[18049] = 16'h495e;
mem_array[18048] = 16'h3e8a;
mem_array[18051] = 16'h0757;
mem_array[18050] = 16'h3e20;
mem_array[18053] = 16'h2864;
mem_array[18052] = 16'hbef1;
mem_array[18055] = 16'h378e;
mem_array[18054] = 16'h3ed3;
mem_array[18057] = 16'h5723;
mem_array[18056] = 16'h3e18;
mem_array[18059] = 16'h43ce;
mem_array[18058] = 16'hbebd;
mem_array[18061] = 16'h7ccd;
mem_array[18060] = 16'h3ed7;
mem_array[18063] = 16'h26c2;
mem_array[18062] = 16'h3e76;
mem_array[18065] = 16'ha3fb;
mem_array[18064] = 16'hbe98;
mem_array[18067] = 16'h5403;
mem_array[18066] = 16'h3e9c;
mem_array[18069] = 16'hb1ef;
mem_array[18068] = 16'hbe39;
mem_array[18071] = 16'h4cd5;
mem_array[18070] = 16'hbf18;
mem_array[18073] = 16'hdb25;
mem_array[18072] = 16'hbebe;
mem_array[18075] = 16'hcbe2;
mem_array[18074] = 16'h3e58;
mem_array[18077] = 16'h89fb;
mem_array[18076] = 16'h3d10;
mem_array[18079] = 16'h5cce;
mem_array[18078] = 16'hbe85;
mem_array[18081] = 16'h375e;
mem_array[18080] = 16'h3add;
mem_array[18083] = 16'hb75a;
mem_array[18082] = 16'hbcb4;
mem_array[18085] = 16'h39e6;
mem_array[18084] = 16'hbd34;
mem_array[18087] = 16'h4f77;
mem_array[18086] = 16'hbe01;
mem_array[18089] = 16'ha0c8;
mem_array[18088] = 16'h3ec0;
mem_array[18091] = 16'h17f8;
mem_array[18090] = 16'h3da2;
mem_array[18093] = 16'hecf1;
mem_array[18092] = 16'h3e44;
mem_array[18095] = 16'hd773;
mem_array[18094] = 16'hbe5f;
mem_array[18097] = 16'hced5;
mem_array[18096] = 16'hbe84;
mem_array[18099] = 16'h7db6;
mem_array[18098] = 16'h3df7;
mem_array[18101] = 16'h7d44;
mem_array[18100] = 16'hbe02;
mem_array[18103] = 16'h6245;
mem_array[18102] = 16'hbd75;
mem_array[18105] = 16'hbcdb;
mem_array[18104] = 16'hbfbc;
mem_array[18107] = 16'hccc3;
mem_array[18106] = 16'hbd27;
mem_array[18109] = 16'h7599;
mem_array[18108] = 16'h3e83;
mem_array[18111] = 16'h6e8f;
mem_array[18110] = 16'h3d97;
mem_array[18113] = 16'h4e48;
mem_array[18112] = 16'hbea3;
mem_array[18115] = 16'h0653;
mem_array[18114] = 16'h3f17;
mem_array[18117] = 16'he0d1;
mem_array[18116] = 16'hbd55;
mem_array[18119] = 16'h88dd;
mem_array[18118] = 16'hbf1d;
mem_array[18121] = 16'h9664;
mem_array[18120] = 16'h3e17;
mem_array[18123] = 16'hcec0;
mem_array[18122] = 16'h3ec3;
mem_array[18125] = 16'h9155;
mem_array[18124] = 16'hbe54;
mem_array[18127] = 16'h151f;
mem_array[18126] = 16'h3f0d;
mem_array[18129] = 16'h7468;
mem_array[18128] = 16'hbe45;
mem_array[18131] = 16'h15cb;
mem_array[18130] = 16'hbe90;
mem_array[18133] = 16'hb51f;
mem_array[18132] = 16'hbe89;
mem_array[18135] = 16'h2799;
mem_array[18134] = 16'h3e54;
mem_array[18137] = 16'h0856;
mem_array[18136] = 16'h3d5c;
mem_array[18139] = 16'hcf27;
mem_array[18138] = 16'h3f6b;
mem_array[18141] = 16'hedda;
mem_array[18140] = 16'hbc88;
mem_array[18143] = 16'h3c17;
mem_array[18142] = 16'hbd4d;
mem_array[18145] = 16'hc6c2;
mem_array[18144] = 16'hbe65;
mem_array[18147] = 16'hbd63;
mem_array[18146] = 16'hbd77;
mem_array[18149] = 16'h1f7f;
mem_array[18148] = 16'hbe97;
mem_array[18151] = 16'h4a31;
mem_array[18150] = 16'h3ee7;
mem_array[18153] = 16'h7772;
mem_array[18152] = 16'hbef3;
mem_array[18155] = 16'he29b;
mem_array[18154] = 16'hbe33;
mem_array[18157] = 16'h2a05;
mem_array[18156] = 16'hbc74;
mem_array[18159] = 16'hddf7;
mem_array[18158] = 16'hbe63;
mem_array[18161] = 16'h2e88;
mem_array[18160] = 16'hbd51;
mem_array[18163] = 16'h8d5e;
mem_array[18162] = 16'hbe8a;
mem_array[18165] = 16'hc04c;
mem_array[18164] = 16'hbf95;
mem_array[18167] = 16'h237d;
mem_array[18166] = 16'hbe04;
mem_array[18169] = 16'hf3bd;
mem_array[18168] = 16'hbe58;
mem_array[18171] = 16'h2c62;
mem_array[18170] = 16'h3d7a;
mem_array[18173] = 16'he1cb;
mem_array[18172] = 16'hbf12;
mem_array[18175] = 16'he709;
mem_array[18174] = 16'h3f33;
mem_array[18177] = 16'ha2e0;
mem_array[18176] = 16'hbdce;
mem_array[18179] = 16'hd67a;
mem_array[18178] = 16'hbf28;
mem_array[18181] = 16'h1009;
mem_array[18180] = 16'hbf4b;
mem_array[18183] = 16'h4bb1;
mem_array[18182] = 16'h3ef6;
mem_array[18185] = 16'h3e70;
mem_array[18184] = 16'hbe0e;
mem_array[18187] = 16'heae6;
mem_array[18186] = 16'h3f43;
mem_array[18189] = 16'h765b;
mem_array[18188] = 16'h3d9a;
mem_array[18191] = 16'hde3e;
mem_array[18190] = 16'hbf19;
mem_array[18193] = 16'h3885;
mem_array[18192] = 16'hbfc3;
mem_array[18195] = 16'hb83d;
mem_array[18194] = 16'hbe3a;
mem_array[18197] = 16'h6199;
mem_array[18196] = 16'hbe10;
mem_array[18199] = 16'h4c67;
mem_array[18198] = 16'hbe6d;
mem_array[18201] = 16'h56b7;
mem_array[18200] = 16'h3d68;
mem_array[18203] = 16'h3d91;
mem_array[18202] = 16'hbc9b;
mem_array[18205] = 16'hcf87;
mem_array[18204] = 16'hbed8;
mem_array[18207] = 16'h6d53;
mem_array[18206] = 16'hbf69;
mem_array[18209] = 16'h135f;
mem_array[18208] = 16'h3e2f;
mem_array[18211] = 16'h16e4;
mem_array[18210] = 16'h3e84;
mem_array[18213] = 16'heb7e;
mem_array[18212] = 16'hbf26;
mem_array[18215] = 16'h5364;
mem_array[18214] = 16'hbf06;
mem_array[18217] = 16'h021c;
mem_array[18216] = 16'hbed0;
mem_array[18219] = 16'h5bca;
mem_array[18218] = 16'hbee4;
mem_array[18221] = 16'h5307;
mem_array[18220] = 16'hbdd3;
mem_array[18223] = 16'hf19b;
mem_array[18222] = 16'hbdfe;
mem_array[18225] = 16'h7682;
mem_array[18224] = 16'hbf64;
mem_array[18227] = 16'heccb;
mem_array[18226] = 16'h3e6e;
mem_array[18229] = 16'h1954;
mem_array[18228] = 16'hbf26;
mem_array[18231] = 16'h63e5;
mem_array[18230] = 16'hbea5;
mem_array[18233] = 16'h3fc9;
mem_array[18232] = 16'h3e31;
mem_array[18235] = 16'hced6;
mem_array[18234] = 16'h3f4c;
mem_array[18237] = 16'h2173;
mem_array[18236] = 16'hbfad;
mem_array[18239] = 16'h4ecb;
mem_array[18238] = 16'hbfa9;
mem_array[18241] = 16'h6839;
mem_array[18240] = 16'hc017;
mem_array[18243] = 16'hec51;
mem_array[18242] = 16'hbe90;
mem_array[18245] = 16'h7a93;
mem_array[18244] = 16'h3eec;
mem_array[18247] = 16'h2acc;
mem_array[18246] = 16'hbd80;
mem_array[18249] = 16'h0d17;
mem_array[18248] = 16'h3dee;
mem_array[18251] = 16'hf8ae;
mem_array[18250] = 16'h3d99;
mem_array[18253] = 16'h1c87;
mem_array[18252] = 16'hbfcc;
mem_array[18255] = 16'h4fb9;
mem_array[18254] = 16'h3ea2;
mem_array[18257] = 16'hf066;
mem_array[18256] = 16'hbebf;
mem_array[18259] = 16'he128;
mem_array[18258] = 16'hbf02;
mem_array[18261] = 16'h0adc;
mem_array[18260] = 16'hbdf4;
mem_array[18263] = 16'h576a;
mem_array[18262] = 16'h3987;
mem_array[18265] = 16'hb69f;
mem_array[18264] = 16'hbf82;
mem_array[18267] = 16'h60c3;
mem_array[18266] = 16'hbf23;
mem_array[18269] = 16'hc212;
mem_array[18268] = 16'h3f47;
mem_array[18271] = 16'hb889;
mem_array[18270] = 16'hbeb6;
mem_array[18273] = 16'he118;
mem_array[18272] = 16'hbf10;
mem_array[18275] = 16'h2a47;
mem_array[18274] = 16'h3f00;
mem_array[18277] = 16'h6eff;
mem_array[18276] = 16'hbecb;
mem_array[18279] = 16'h16ba;
mem_array[18278] = 16'h3ec9;
mem_array[18281] = 16'h7e87;
mem_array[18280] = 16'hbf09;
mem_array[18283] = 16'h5535;
mem_array[18282] = 16'h3eb2;
mem_array[18285] = 16'h0d02;
mem_array[18284] = 16'hbf02;
mem_array[18287] = 16'h247f;
mem_array[18286] = 16'hbe48;
mem_array[18289] = 16'had98;
mem_array[18288] = 16'hbf19;
mem_array[18291] = 16'hf643;
mem_array[18290] = 16'h3e8a;
mem_array[18293] = 16'h2fe3;
mem_array[18292] = 16'h3c9a;
mem_array[18295] = 16'h4a75;
mem_array[18294] = 16'h3f81;
mem_array[18297] = 16'h8369;
mem_array[18296] = 16'hbf81;
mem_array[18299] = 16'h9cd3;
mem_array[18298] = 16'hbfb1;
mem_array[18301] = 16'h7d38;
mem_array[18300] = 16'hbf92;
mem_array[18303] = 16'h084b;
mem_array[18302] = 16'h3e9f;
mem_array[18305] = 16'h74c3;
mem_array[18304] = 16'hbe8d;
mem_array[18307] = 16'hed51;
mem_array[18306] = 16'hbf99;
mem_array[18309] = 16'h8701;
mem_array[18308] = 16'h3e86;
mem_array[18311] = 16'h20e1;
mem_array[18310] = 16'h3e98;
mem_array[18313] = 16'h4eb4;
mem_array[18312] = 16'hbef7;
mem_array[18315] = 16'h6118;
mem_array[18314] = 16'h3f12;
mem_array[18317] = 16'h3d2b;
mem_array[18316] = 16'hbeb1;
mem_array[18319] = 16'h6651;
mem_array[18318] = 16'h3f21;
mem_array[18321] = 16'haf0c;
mem_array[18320] = 16'hbcf4;
mem_array[18323] = 16'h8050;
mem_array[18322] = 16'h3d80;
mem_array[18325] = 16'h34f1;
mem_array[18324] = 16'hbf5e;
mem_array[18327] = 16'hceed;
mem_array[18326] = 16'hbe89;
mem_array[18329] = 16'h8871;
mem_array[18328] = 16'hbf07;
mem_array[18331] = 16'hc58c;
mem_array[18330] = 16'hbe12;
mem_array[18333] = 16'hc3f9;
mem_array[18332] = 16'hbee2;
mem_array[18335] = 16'h5419;
mem_array[18334] = 16'h3f52;
mem_array[18337] = 16'h73bc;
mem_array[18336] = 16'h3eda;
mem_array[18339] = 16'hbfef;
mem_array[18338] = 16'h3da0;
mem_array[18341] = 16'hf54e;
mem_array[18340] = 16'h3ed3;
mem_array[18343] = 16'ha905;
mem_array[18342] = 16'h3eaa;
mem_array[18345] = 16'h9d07;
mem_array[18344] = 16'hbf4a;
mem_array[18347] = 16'h6617;
mem_array[18346] = 16'hbf12;
mem_array[18349] = 16'h44f2;
mem_array[18348] = 16'h3b83;
mem_array[18351] = 16'h0b57;
mem_array[18350] = 16'h3c21;
mem_array[18353] = 16'h8a1c;
mem_array[18352] = 16'hbda8;
mem_array[18355] = 16'h9872;
mem_array[18354] = 16'h3f79;
mem_array[18357] = 16'h11df;
mem_array[18356] = 16'hbf23;
mem_array[18359] = 16'hc67a;
mem_array[18358] = 16'hbf7d;
mem_array[18361] = 16'hf88e;
mem_array[18360] = 16'h3f1b;
mem_array[18363] = 16'h58b6;
mem_array[18362] = 16'hbf2a;
mem_array[18365] = 16'hca5a;
mem_array[18364] = 16'h3ebd;
mem_array[18367] = 16'hf3af;
mem_array[18366] = 16'hbf9f;
mem_array[18369] = 16'h43b2;
mem_array[18368] = 16'hbfb0;
mem_array[18371] = 16'h8208;
mem_array[18370] = 16'h3f4c;
mem_array[18373] = 16'h75b3;
mem_array[18372] = 16'h3e1d;
mem_array[18375] = 16'h9d0e;
mem_array[18374] = 16'hbebb;
mem_array[18377] = 16'h651c;
mem_array[18376] = 16'hbe66;
mem_array[18379] = 16'h1ea7;
mem_array[18378] = 16'hbd9f;
mem_array[18381] = 16'haba8;
mem_array[18380] = 16'hbbf3;
mem_array[18383] = 16'h2d5c;
mem_array[18382] = 16'hbcd8;
mem_array[18385] = 16'h8c41;
mem_array[18384] = 16'hbf22;
mem_array[18387] = 16'h9504;
mem_array[18386] = 16'h3db7;
mem_array[18389] = 16'h12f6;
mem_array[18388] = 16'h3ec6;
mem_array[18391] = 16'h866b;
mem_array[18390] = 16'hbe48;
mem_array[18393] = 16'h3a6a;
mem_array[18392] = 16'hbe8a;
mem_array[18395] = 16'hc545;
mem_array[18394] = 16'hbecb;
mem_array[18397] = 16'h3d79;
mem_array[18396] = 16'hbf54;
mem_array[18399] = 16'h446b;
mem_array[18398] = 16'hbda8;
mem_array[18401] = 16'h1a92;
mem_array[18400] = 16'hc003;
mem_array[18403] = 16'hbd06;
mem_array[18402] = 16'hbdc2;
mem_array[18405] = 16'h9023;
mem_array[18404] = 16'h3e31;
mem_array[18407] = 16'h10e0;
mem_array[18406] = 16'hbee0;
mem_array[18409] = 16'h1f30;
mem_array[18408] = 16'h3eca;
mem_array[18411] = 16'h71c3;
mem_array[18410] = 16'hbee5;
mem_array[18413] = 16'h4e16;
mem_array[18412] = 16'h3f69;
mem_array[18415] = 16'h3534;
mem_array[18414] = 16'h3ee5;
mem_array[18417] = 16'h80ee;
mem_array[18416] = 16'h3ea2;
mem_array[18419] = 16'hf1e8;
mem_array[18418] = 16'hbfa4;
mem_array[18421] = 16'h5c20;
mem_array[18420] = 16'h3f31;
mem_array[18423] = 16'h33ba;
mem_array[18422] = 16'hbef0;
mem_array[18425] = 16'hc178;
mem_array[18424] = 16'hbe05;
mem_array[18427] = 16'hc4fd;
mem_array[18426] = 16'hbdad;
mem_array[18429] = 16'h5a68;
mem_array[18428] = 16'h3d46;
mem_array[18431] = 16'h06f7;
mem_array[18430] = 16'h3f88;
mem_array[18433] = 16'h9cf0;
mem_array[18432] = 16'hbe0b;
mem_array[18435] = 16'h4d4a;
mem_array[18434] = 16'h3d14;
mem_array[18437] = 16'h1675;
mem_array[18436] = 16'h3df2;
mem_array[18439] = 16'h51c6;
mem_array[18438] = 16'h3f18;
mem_array[18441] = 16'h4bcc;
mem_array[18440] = 16'hbd7e;
mem_array[18443] = 16'ha0f1;
mem_array[18442] = 16'hbca3;
mem_array[18445] = 16'h4642;
mem_array[18444] = 16'hbe5d;
mem_array[18447] = 16'h39c0;
mem_array[18446] = 16'h3d6d;
mem_array[18449] = 16'h03fb;
mem_array[18448] = 16'hbbb5;
mem_array[18451] = 16'h4072;
mem_array[18450] = 16'h3e89;
mem_array[18453] = 16'ha180;
mem_array[18452] = 16'hbc6b;
mem_array[18455] = 16'hd66c;
mem_array[18454] = 16'h3e2b;
mem_array[18457] = 16'h1637;
mem_array[18456] = 16'hbe43;
mem_array[18459] = 16'h9ad2;
mem_array[18458] = 16'hbdad;
mem_array[18461] = 16'h208d;
mem_array[18460] = 16'hbe58;
mem_array[18463] = 16'h15c6;
mem_array[18462] = 16'h3e04;
mem_array[18465] = 16'hefe8;
mem_array[18464] = 16'hbd3a;
mem_array[18467] = 16'h1c9d;
mem_array[18466] = 16'hbf19;
mem_array[18469] = 16'hd0ac;
mem_array[18468] = 16'hbdf5;
mem_array[18471] = 16'h45f5;
mem_array[18470] = 16'hbd49;
mem_array[18473] = 16'h5b2a;
mem_array[18472] = 16'h3eb0;
mem_array[18475] = 16'hf9a5;
mem_array[18474] = 16'h3f05;
mem_array[18477] = 16'h01cc;
mem_array[18476] = 16'h3d36;
mem_array[18479] = 16'h837d;
mem_array[18478] = 16'hbedd;
mem_array[18481] = 16'he9b0;
mem_array[18480] = 16'h3d4a;
mem_array[18483] = 16'h3d0f;
mem_array[18482] = 16'hbb8b;
mem_array[18485] = 16'h634b;
mem_array[18484] = 16'h3d25;
mem_array[18487] = 16'hc3b5;
mem_array[18486] = 16'h3da4;
mem_array[18489] = 16'hbec5;
mem_array[18488] = 16'h3d13;
mem_array[18491] = 16'h9434;
mem_array[18490] = 16'hbb26;
mem_array[18493] = 16'hddec;
mem_array[18492] = 16'hbdbc;
mem_array[18495] = 16'h5163;
mem_array[18494] = 16'hbda5;
mem_array[18497] = 16'h4099;
mem_array[18496] = 16'h3d59;
mem_array[18499] = 16'h0feb;
mem_array[18498] = 16'hbc51;
mem_array[18501] = 16'h4627;
mem_array[18500] = 16'hbca3;
mem_array[18503] = 16'h8dd0;
mem_array[18502] = 16'h3da2;
mem_array[18505] = 16'hccf0;
mem_array[18504] = 16'h3d6b;
mem_array[18507] = 16'h9b93;
mem_array[18506] = 16'hbd1b;
mem_array[18509] = 16'ha9b1;
mem_array[18508] = 16'hbd53;
mem_array[18511] = 16'ha569;
mem_array[18510] = 16'hbd97;
mem_array[18513] = 16'h1cec;
mem_array[18512] = 16'hbd3a;
mem_array[18515] = 16'hbcda;
mem_array[18514] = 16'hbcbb;
mem_array[18517] = 16'hd853;
mem_array[18516] = 16'h3e1c;
mem_array[18519] = 16'h5eaa;
mem_array[18518] = 16'h3e45;
mem_array[18521] = 16'he3c0;
mem_array[18520] = 16'hbda0;
mem_array[18523] = 16'h34eb;
mem_array[18522] = 16'h3cd2;
mem_array[18525] = 16'h157c;
mem_array[18524] = 16'hbd32;
mem_array[18527] = 16'h4537;
mem_array[18526] = 16'hbde1;
mem_array[18529] = 16'h70de;
mem_array[18528] = 16'hbd1f;
mem_array[18531] = 16'hd4da;
mem_array[18530] = 16'h3d28;
mem_array[18533] = 16'h0276;
mem_array[18532] = 16'hbe1a;
mem_array[18535] = 16'hc3cf;
mem_array[18534] = 16'h3e28;
mem_array[18537] = 16'h1040;
mem_array[18536] = 16'hbd8d;
mem_array[18539] = 16'hdf06;
mem_array[18538] = 16'hbdbe;
mem_array[18541] = 16'hf6fc;
mem_array[18540] = 16'h3e27;
mem_array[18543] = 16'h3a69;
mem_array[18542] = 16'h3f43;
mem_array[18545] = 16'he4d9;
mem_array[18544] = 16'h3e8d;
mem_array[18547] = 16'hebdb;
mem_array[18546] = 16'h3ec4;
mem_array[18549] = 16'he5f5;
mem_array[18548] = 16'hbf16;
mem_array[18551] = 16'hb886;
mem_array[18550] = 16'hbe1f;
mem_array[18553] = 16'h4c58;
mem_array[18552] = 16'hbd38;
mem_array[18555] = 16'h599f;
mem_array[18554] = 16'h3dc6;
mem_array[18557] = 16'h6c32;
mem_array[18556] = 16'hbe51;
mem_array[18559] = 16'h76c2;
mem_array[18558] = 16'h3e59;
mem_array[18561] = 16'h7923;
mem_array[18560] = 16'h39a3;
mem_array[18563] = 16'h96c1;
mem_array[18562] = 16'hbcd1;
mem_array[18565] = 16'h8b59;
mem_array[18564] = 16'h3f46;
mem_array[18567] = 16'h2e4e;
mem_array[18566] = 16'hbded;
mem_array[18569] = 16'h54a8;
mem_array[18568] = 16'hbd75;
mem_array[18571] = 16'h3686;
mem_array[18570] = 16'hbf3d;
mem_array[18573] = 16'hffce;
mem_array[18572] = 16'h3e58;
mem_array[18575] = 16'h85bc;
mem_array[18574] = 16'hbeb0;
mem_array[18577] = 16'hb9da;
mem_array[18576] = 16'hbe68;
mem_array[18579] = 16'hcba1;
mem_array[18578] = 16'h3d74;
mem_array[18581] = 16'he697;
mem_array[18580] = 16'hbdd0;
mem_array[18583] = 16'h69ae;
mem_array[18582] = 16'h3f12;
mem_array[18585] = 16'hfc45;
mem_array[18584] = 16'hbccf;
mem_array[18587] = 16'h5e93;
mem_array[18586] = 16'h3ebc;
mem_array[18589] = 16'h08b2;
mem_array[18588] = 16'hbe69;
mem_array[18591] = 16'hd9fa;
mem_array[18590] = 16'h3f89;
mem_array[18593] = 16'h6f44;
mem_array[18592] = 16'hbe81;
mem_array[18595] = 16'h1298;
mem_array[18594] = 16'h3ead;
mem_array[18597] = 16'hcc61;
mem_array[18596] = 16'h3d12;
mem_array[18599] = 16'h9f02;
mem_array[18598] = 16'hbe91;
mem_array[18601] = 16'h1bd1;
mem_array[18600] = 16'h3e1c;
mem_array[18603] = 16'hc1e2;
mem_array[18602] = 16'h3ef6;
mem_array[18605] = 16'h4124;
mem_array[18604] = 16'hbe44;
mem_array[18607] = 16'hc5e2;
mem_array[18606] = 16'h3da0;
mem_array[18609] = 16'hfe94;
mem_array[18608] = 16'h3e04;
mem_array[18611] = 16'h84b2;
mem_array[18610] = 16'h3e5c;
mem_array[18613] = 16'h8050;
mem_array[18612] = 16'hbed2;
mem_array[18615] = 16'h070e;
mem_array[18614] = 16'hbd79;
mem_array[18617] = 16'h87f4;
mem_array[18616] = 16'hbf2a;
mem_array[18619] = 16'h54a6;
mem_array[18618] = 16'h3f1a;
mem_array[18621] = 16'hf304;
mem_array[18620] = 16'hbde7;
mem_array[18623] = 16'hc9ab;
mem_array[18622] = 16'hbd1f;
mem_array[18625] = 16'hc5f7;
mem_array[18624] = 16'h3ec3;
mem_array[18627] = 16'ha30e;
mem_array[18626] = 16'hbf0a;
mem_array[18629] = 16'hb590;
mem_array[18628] = 16'hbf16;
mem_array[18631] = 16'h97de;
mem_array[18630] = 16'hbd78;
mem_array[18633] = 16'hf964;
mem_array[18632] = 16'hbe90;
mem_array[18635] = 16'h7b57;
mem_array[18634] = 16'hbed8;
mem_array[18637] = 16'h782f;
mem_array[18636] = 16'h3f0e;
mem_array[18639] = 16'hcf72;
mem_array[18638] = 16'hbead;
mem_array[18641] = 16'h5832;
mem_array[18640] = 16'hbf29;
mem_array[18643] = 16'h18fe;
mem_array[18642] = 16'h3dd1;
mem_array[18645] = 16'h8e84;
mem_array[18644] = 16'h3ce9;
mem_array[18647] = 16'h2e52;
mem_array[18646] = 16'h3f12;
mem_array[18649] = 16'ha8d0;
mem_array[18648] = 16'hbf8a;
mem_array[18651] = 16'hb980;
mem_array[18650] = 16'h3f0e;
mem_array[18653] = 16'hf934;
mem_array[18652] = 16'hbeec;
mem_array[18655] = 16'haa4d;
mem_array[18654] = 16'h3ec8;
mem_array[18657] = 16'h918a;
mem_array[18656] = 16'hbf15;
mem_array[18659] = 16'h6df6;
mem_array[18658] = 16'hbf06;
mem_array[18661] = 16'h7106;
mem_array[18660] = 16'hbe8c;
mem_array[18663] = 16'h95e0;
mem_array[18662] = 16'h3f5b;
mem_array[18665] = 16'h93d2;
mem_array[18664] = 16'h3dd6;
mem_array[18667] = 16'h4779;
mem_array[18666] = 16'hbf85;
mem_array[18669] = 16'h5d4f;
mem_array[18668] = 16'hbde9;
mem_array[18671] = 16'hdea1;
mem_array[18670] = 16'h3f3a;
mem_array[18673] = 16'h2fce;
mem_array[18672] = 16'hbf73;
mem_array[18675] = 16'hf8e2;
mem_array[18674] = 16'h3e90;
mem_array[18677] = 16'he368;
mem_array[18676] = 16'h3e89;
mem_array[18679] = 16'h2b19;
mem_array[18678] = 16'hbf19;
mem_array[18681] = 16'hfd12;
mem_array[18680] = 16'hbc79;
mem_array[18683] = 16'h0e75;
mem_array[18682] = 16'h3cd7;
mem_array[18685] = 16'h1b9b;
mem_array[18684] = 16'hbf6a;
mem_array[18687] = 16'haf39;
mem_array[18686] = 16'hbeca;
mem_array[18689] = 16'h3478;
mem_array[18688] = 16'h3dc4;
mem_array[18691] = 16'h76d8;
mem_array[18690] = 16'h3ea4;
mem_array[18693] = 16'h93dc;
mem_array[18692] = 16'h3e7c;
mem_array[18695] = 16'hc9f8;
mem_array[18694] = 16'h3ee8;
mem_array[18697] = 16'hf75e;
mem_array[18696] = 16'h3f33;
mem_array[18699] = 16'h65e2;
mem_array[18698] = 16'hbe6c;
mem_array[18701] = 16'h3315;
mem_array[18700] = 16'hbf7e;
mem_array[18703] = 16'heaa9;
mem_array[18702] = 16'hbe18;
mem_array[18705] = 16'h25eb;
mem_array[18704] = 16'hbf5d;
mem_array[18707] = 16'h12ad;
mem_array[18706] = 16'hbe5b;
mem_array[18709] = 16'h46af;
mem_array[18708] = 16'h3e39;
mem_array[18711] = 16'h17bc;
mem_array[18710] = 16'h3e11;
mem_array[18713] = 16'h1244;
mem_array[18712] = 16'h3e1a;
mem_array[18715] = 16'h4400;
mem_array[18714] = 16'h3e41;
mem_array[18717] = 16'habf8;
mem_array[18716] = 16'hbf1f;
mem_array[18719] = 16'h9d48;
mem_array[18718] = 16'h3e62;
mem_array[18721] = 16'h31c7;
mem_array[18720] = 16'h3f2d;
mem_array[18723] = 16'hf153;
mem_array[18722] = 16'h3e10;
mem_array[18725] = 16'h6929;
mem_array[18724] = 16'h3f14;
mem_array[18727] = 16'h6dce;
mem_array[18726] = 16'hbdcf;
mem_array[18729] = 16'h3983;
mem_array[18728] = 16'hbed7;
mem_array[18731] = 16'h5bd8;
mem_array[18730] = 16'h3f0e;
mem_array[18733] = 16'h9bf8;
mem_array[18732] = 16'hbf97;
mem_array[18735] = 16'h9c6f;
mem_array[18734] = 16'h3e14;
mem_array[18737] = 16'h3744;
mem_array[18736] = 16'hbf57;
mem_array[18739] = 16'he356;
mem_array[18738] = 16'hbd5f;
mem_array[18741] = 16'h3d0e;
mem_array[18740] = 16'hbd28;
mem_array[18743] = 16'h873f;
mem_array[18742] = 16'h39eb;
mem_array[18745] = 16'h622a;
mem_array[18744] = 16'hbf18;
mem_array[18747] = 16'hf784;
mem_array[18746] = 16'hbec3;
mem_array[18749] = 16'h11a3;
mem_array[18748] = 16'h3dc5;
mem_array[18751] = 16'h1fd9;
mem_array[18750] = 16'hbe67;
mem_array[18753] = 16'he5a9;
mem_array[18752] = 16'h3f90;
mem_array[18755] = 16'h42b8;
mem_array[18754] = 16'hbdcd;
mem_array[18757] = 16'hb164;
mem_array[18756] = 16'h3e2c;
mem_array[18759] = 16'h8c47;
mem_array[18758] = 16'hbe20;
mem_array[18761] = 16'hb667;
mem_array[18760] = 16'hbef4;
mem_array[18763] = 16'h5cc4;
mem_array[18762] = 16'h3e37;
mem_array[18765] = 16'h314c;
mem_array[18764] = 16'hbf17;
mem_array[18767] = 16'h7b9f;
mem_array[18766] = 16'h3d66;
mem_array[18769] = 16'h1f92;
mem_array[18768] = 16'h3f37;
mem_array[18771] = 16'haa5d;
mem_array[18770] = 16'h3ee1;
mem_array[18773] = 16'hbe04;
mem_array[18772] = 16'h3f21;
mem_array[18775] = 16'hdd4d;
mem_array[18774] = 16'hbe83;
mem_array[18777] = 16'hf682;
mem_array[18776] = 16'hbf5d;
mem_array[18779] = 16'ha75c;
mem_array[18778] = 16'hbeae;
mem_array[18781] = 16'h2161;
mem_array[18780] = 16'hbb01;
mem_array[18783] = 16'h160c;
mem_array[18782] = 16'h3dfa;
mem_array[18785] = 16'hf6a1;
mem_array[18784] = 16'h3e05;
mem_array[18787] = 16'h7ee3;
mem_array[18786] = 16'hbf19;
mem_array[18789] = 16'h32df;
mem_array[18788] = 16'hbe47;
mem_array[18791] = 16'h610b;
mem_array[18790] = 16'hbe0d;
mem_array[18793] = 16'h89fb;
mem_array[18792] = 16'hbfe6;
mem_array[18795] = 16'h3ae7;
mem_array[18794] = 16'hbe59;
mem_array[18797] = 16'hfe35;
mem_array[18796] = 16'h3ee4;
mem_array[18799] = 16'h199f;
mem_array[18798] = 16'h3ecc;
mem_array[18801] = 16'he0c7;
mem_array[18800] = 16'h3c9c;
mem_array[18803] = 16'h23c7;
mem_array[18802] = 16'h3bca;
mem_array[18805] = 16'h2fd4;
mem_array[18804] = 16'hbec3;
mem_array[18807] = 16'h2851;
mem_array[18806] = 16'hbe9a;
mem_array[18809] = 16'ha879;
mem_array[18808] = 16'h3de7;
mem_array[18811] = 16'hf6f7;
mem_array[18810] = 16'h3ead;
mem_array[18813] = 16'h4268;
mem_array[18812] = 16'h3f37;
mem_array[18815] = 16'h019c;
mem_array[18814] = 16'h3e54;
mem_array[18817] = 16'h25c8;
mem_array[18816] = 16'h3e5d;
mem_array[18819] = 16'h8b02;
mem_array[18818] = 16'h3d2e;
mem_array[18821] = 16'ha297;
mem_array[18820] = 16'hbe31;
mem_array[18823] = 16'h234f;
mem_array[18822] = 16'hbdf6;
mem_array[18825] = 16'hd4c8;
mem_array[18824] = 16'hbea9;
mem_array[18827] = 16'hb0a6;
mem_array[18826] = 16'hbe6a;
mem_array[18829] = 16'h49f1;
mem_array[18828] = 16'hba9d;
mem_array[18831] = 16'h8965;
mem_array[18830] = 16'h3dab;
mem_array[18833] = 16'hb481;
mem_array[18832] = 16'hbde4;
mem_array[18835] = 16'hcd6d;
mem_array[18834] = 16'hbee9;
mem_array[18837] = 16'h507e;
mem_array[18836] = 16'hbf46;
mem_array[18839] = 16'h0df9;
mem_array[18838] = 16'h3df0;
mem_array[18841] = 16'hf8ae;
mem_array[18840] = 16'hbe90;
mem_array[18843] = 16'h5a1e;
mem_array[18842] = 16'h3c8c;
mem_array[18845] = 16'hf1f6;
mem_array[18844] = 16'h3ec8;
mem_array[18847] = 16'h31dd;
mem_array[18846] = 16'hbf00;
mem_array[18849] = 16'ha898;
mem_array[18848] = 16'h3d5f;
mem_array[18851] = 16'h14eb;
mem_array[18850] = 16'hbcc9;
mem_array[18853] = 16'h5de8;
mem_array[18852] = 16'hbfc8;
mem_array[18855] = 16'h68e5;
mem_array[18854] = 16'hbe75;
mem_array[18857] = 16'hfef4;
mem_array[18856] = 16'hbd82;
mem_array[18859] = 16'h843f;
mem_array[18858] = 16'h3d10;
mem_array[18861] = 16'he888;
mem_array[18860] = 16'hbd82;
mem_array[18863] = 16'hf5c8;
mem_array[18862] = 16'hbdab;
mem_array[18865] = 16'he1f8;
mem_array[18864] = 16'hbdd2;
mem_array[18867] = 16'hc677;
mem_array[18866] = 16'hbf6c;
mem_array[18869] = 16'h670d;
mem_array[18868] = 16'hbe38;
mem_array[18871] = 16'had04;
mem_array[18870] = 16'h3dce;
mem_array[18873] = 16'hf99e;
mem_array[18872] = 16'h3f15;
mem_array[18875] = 16'h8cde;
mem_array[18874] = 16'h3d9a;
mem_array[18877] = 16'h6d01;
mem_array[18876] = 16'h3e0d;
mem_array[18879] = 16'h37aa;
mem_array[18878] = 16'h3dda;
mem_array[18881] = 16'h10c0;
mem_array[18880] = 16'h3e0a;
mem_array[18883] = 16'hda62;
mem_array[18882] = 16'h3e0a;
mem_array[18885] = 16'h356b;
mem_array[18884] = 16'hbecb;
mem_array[18887] = 16'h5b09;
mem_array[18886] = 16'h3e7b;
mem_array[18889] = 16'h3a3e;
mem_array[18888] = 16'h3f39;
mem_array[18891] = 16'h45df;
mem_array[18890] = 16'h3e92;
mem_array[18893] = 16'ha4ad;
mem_array[18892] = 16'h3e28;
mem_array[18895] = 16'h9917;
mem_array[18894] = 16'hbe7f;
mem_array[18897] = 16'hd1a6;
mem_array[18896] = 16'hbf6b;
mem_array[18899] = 16'h131b;
mem_array[18898] = 16'h3d05;
mem_array[18901] = 16'hf947;
mem_array[18900] = 16'hbf28;
mem_array[18903] = 16'h3c44;
mem_array[18902] = 16'h3d0b;
mem_array[18905] = 16'hd5c9;
mem_array[18904] = 16'h3e90;
mem_array[18907] = 16'h085e;
mem_array[18906] = 16'h3d3e;
mem_array[18909] = 16'h371c;
mem_array[18908] = 16'hbe16;
mem_array[18911] = 16'h7b15;
mem_array[18910] = 16'h3ed4;
mem_array[18913] = 16'h65f9;
mem_array[18912] = 16'hbfcf;
mem_array[18915] = 16'h0306;
mem_array[18914] = 16'h3f04;
mem_array[18917] = 16'h6b6c;
mem_array[18916] = 16'h3ee1;
mem_array[18919] = 16'h00b0;
mem_array[18918] = 16'hbe11;
mem_array[18921] = 16'h69e0;
mem_array[18920] = 16'h3cae;
mem_array[18923] = 16'h545c;
mem_array[18922] = 16'hbd5d;
mem_array[18925] = 16'h4a5c;
mem_array[18924] = 16'hbe51;
mem_array[18927] = 16'h35f3;
mem_array[18926] = 16'hbf4b;
mem_array[18929] = 16'ha034;
mem_array[18928] = 16'hbe17;
mem_array[18931] = 16'hadce;
mem_array[18930] = 16'h3e51;
mem_array[18933] = 16'h6245;
mem_array[18932] = 16'h3e82;
mem_array[18935] = 16'hb0c4;
mem_array[18934] = 16'h3b03;
mem_array[18937] = 16'h42c9;
mem_array[18936] = 16'h3e8d;
mem_array[18939] = 16'hbfe7;
mem_array[18938] = 16'h3c96;
mem_array[18941] = 16'hac34;
mem_array[18940] = 16'hbe1c;
mem_array[18943] = 16'hbe75;
mem_array[18942] = 16'hbd68;
mem_array[18945] = 16'h5d01;
mem_array[18944] = 16'hbf08;
mem_array[18947] = 16'hc3ef;
mem_array[18946] = 16'hbc4c;
mem_array[18949] = 16'hac41;
mem_array[18948] = 16'h3f19;
mem_array[18951] = 16'hd6e7;
mem_array[18950] = 16'hbda4;
mem_array[18953] = 16'h70f2;
mem_array[18952] = 16'hbc8d;
mem_array[18955] = 16'h4675;
mem_array[18954] = 16'hbdcf;
mem_array[18957] = 16'h95a0;
mem_array[18956] = 16'hbfaa;
mem_array[18959] = 16'he4f8;
mem_array[18958] = 16'h3e1e;
mem_array[18961] = 16'h9c99;
mem_array[18960] = 16'hbf01;
mem_array[18963] = 16'h8cf1;
mem_array[18962] = 16'hbe6a;
mem_array[18965] = 16'h7bc5;
mem_array[18964] = 16'h3ed3;
mem_array[18967] = 16'h0bbd;
mem_array[18966] = 16'hbd41;
mem_array[18969] = 16'h2472;
mem_array[18968] = 16'hbcc6;
mem_array[18971] = 16'haf02;
mem_array[18970] = 16'h3ac0;
mem_array[18973] = 16'h4ee2;
mem_array[18972] = 16'hbf9e;
mem_array[18975] = 16'h5b92;
mem_array[18974] = 16'h3f2d;
mem_array[18977] = 16'h4a15;
mem_array[18976] = 16'h3ec9;
mem_array[18979] = 16'h4a5d;
mem_array[18978] = 16'hbe97;
mem_array[18981] = 16'hbe61;
mem_array[18980] = 16'hbd98;
mem_array[18983] = 16'h31a8;
mem_array[18982] = 16'hbd73;
mem_array[18985] = 16'hc643;
mem_array[18984] = 16'hbecf;
mem_array[18987] = 16'h7f81;
mem_array[18986] = 16'hbfa4;
mem_array[18989] = 16'h5b8f;
mem_array[18988] = 16'hbde7;
mem_array[18991] = 16'h9293;
mem_array[18990] = 16'h3e84;
mem_array[18993] = 16'h1719;
mem_array[18992] = 16'hbeac;
mem_array[18995] = 16'h415c;
mem_array[18994] = 16'h3b3b;
mem_array[18997] = 16'hf73a;
mem_array[18996] = 16'h3e6b;
mem_array[18999] = 16'hfa49;
mem_array[18998] = 16'h3e2a;
mem_array[19001] = 16'hee8f;
mem_array[19000] = 16'h3ec1;
mem_array[19003] = 16'h6588;
mem_array[19002] = 16'hbd90;
mem_array[19005] = 16'hb5fb;
mem_array[19004] = 16'hbeb2;
mem_array[19007] = 16'h29c5;
mem_array[19006] = 16'hbe1d;
mem_array[19009] = 16'h97f8;
mem_array[19008] = 16'hbdd4;
mem_array[19011] = 16'h6426;
mem_array[19010] = 16'hbd86;
mem_array[19013] = 16'h9370;
mem_array[19012] = 16'hbd69;
mem_array[19015] = 16'h8c99;
mem_array[19014] = 16'h3d75;
mem_array[19017] = 16'h3fd6;
mem_array[19016] = 16'hbfaf;
mem_array[19019] = 16'h0cfc;
mem_array[19018] = 16'h3e74;
mem_array[19021] = 16'he879;
mem_array[19020] = 16'hbde2;
mem_array[19023] = 16'h025a;
mem_array[19022] = 16'h3e75;
mem_array[19025] = 16'h1574;
mem_array[19024] = 16'h3e33;
mem_array[19027] = 16'h27e3;
mem_array[19026] = 16'hbe82;
mem_array[19029] = 16'h130d;
mem_array[19028] = 16'h3d7f;
mem_array[19031] = 16'hc4ea;
mem_array[19030] = 16'hbeb8;
mem_array[19033] = 16'h434c;
mem_array[19032] = 16'hbf2a;
mem_array[19035] = 16'hf948;
mem_array[19034] = 16'h3e1a;
mem_array[19037] = 16'hff06;
mem_array[19036] = 16'h3ed4;
mem_array[19039] = 16'he0a9;
mem_array[19038] = 16'hbec7;
mem_array[19041] = 16'h2805;
mem_array[19040] = 16'hbc16;
mem_array[19043] = 16'hdbba;
mem_array[19042] = 16'h3cc1;
mem_array[19045] = 16'h3163;
mem_array[19044] = 16'hbe8e;
mem_array[19047] = 16'hbba9;
mem_array[19046] = 16'hbfc2;
mem_array[19049] = 16'h5cda;
mem_array[19048] = 16'h3e81;
mem_array[19051] = 16'h7729;
mem_array[19050] = 16'h3dfd;
mem_array[19053] = 16'h3a44;
mem_array[19052] = 16'hbe08;
mem_array[19055] = 16'hedef;
mem_array[19054] = 16'h3e4b;
mem_array[19057] = 16'h29c7;
mem_array[19056] = 16'h3d8e;
mem_array[19059] = 16'h1140;
mem_array[19058] = 16'h3bd6;
mem_array[19061] = 16'h0207;
mem_array[19060] = 16'h3e09;
mem_array[19063] = 16'hf540;
mem_array[19062] = 16'h3d73;
mem_array[19065] = 16'hca94;
mem_array[19064] = 16'h3e6d;
mem_array[19067] = 16'hc4b0;
mem_array[19066] = 16'hbdb3;
mem_array[19069] = 16'h8007;
mem_array[19068] = 16'hbfac;
mem_array[19071] = 16'h8716;
mem_array[19070] = 16'h3dbd;
mem_array[19073] = 16'h9483;
mem_array[19072] = 16'hbd83;
mem_array[19075] = 16'h3846;
mem_array[19074] = 16'h3d44;
mem_array[19077] = 16'h9186;
mem_array[19076] = 16'hbf82;
mem_array[19079] = 16'h849b;
mem_array[19078] = 16'hbb95;
mem_array[19081] = 16'h3dbe;
mem_array[19080] = 16'hbe6e;
mem_array[19083] = 16'hfb86;
mem_array[19082] = 16'h3ec1;
mem_array[19085] = 16'h8298;
mem_array[19084] = 16'h3eb3;
mem_array[19087] = 16'h9299;
mem_array[19086] = 16'h3d5b;
mem_array[19089] = 16'h060d;
mem_array[19088] = 16'h3df8;
mem_array[19091] = 16'hc8cc;
mem_array[19090] = 16'hbd32;
mem_array[19093] = 16'ha7e6;
mem_array[19092] = 16'hbe72;
mem_array[19095] = 16'h1ee1;
mem_array[19094] = 16'h3e1d;
mem_array[19097] = 16'hb93c;
mem_array[19096] = 16'h3ee3;
mem_array[19099] = 16'h7a93;
mem_array[19098] = 16'hbd5e;
mem_array[19101] = 16'he025;
mem_array[19100] = 16'h3ce7;
mem_array[19103] = 16'hab2a;
mem_array[19102] = 16'hbd5d;
mem_array[19105] = 16'h5387;
mem_array[19104] = 16'h3e7b;
mem_array[19107] = 16'h9f51;
mem_array[19106] = 16'hbf94;
mem_array[19109] = 16'h4405;
mem_array[19108] = 16'h3efb;
mem_array[19111] = 16'h0573;
mem_array[19110] = 16'hbd9d;
mem_array[19113] = 16'hf579;
mem_array[19112] = 16'hbec9;
mem_array[19115] = 16'h591b;
mem_array[19114] = 16'h3eaf;
mem_array[19117] = 16'h9d04;
mem_array[19116] = 16'h3de3;
mem_array[19119] = 16'ha238;
mem_array[19118] = 16'h3e38;
mem_array[19121] = 16'h4ea4;
mem_array[19120] = 16'h3e7f;
mem_array[19123] = 16'h4e95;
mem_array[19122] = 16'hbd9a;
mem_array[19125] = 16'hec7d;
mem_array[19124] = 16'h3d39;
mem_array[19127] = 16'hba44;
mem_array[19126] = 16'hbc39;
mem_array[19129] = 16'h3775;
mem_array[19128] = 16'hc01b;
mem_array[19131] = 16'hda53;
mem_array[19130] = 16'h3e38;
mem_array[19133] = 16'hbee5;
mem_array[19132] = 16'hbddb;
mem_array[19135] = 16'h96d0;
mem_array[19134] = 16'hbaee;
mem_array[19137] = 16'h48cb;
mem_array[19136] = 16'hbf8f;
mem_array[19139] = 16'h15a7;
mem_array[19138] = 16'h3c67;
mem_array[19141] = 16'h4417;
mem_array[19140] = 16'hbef1;
mem_array[19143] = 16'h8b93;
mem_array[19142] = 16'h3eb2;
mem_array[19145] = 16'h3bcf;
mem_array[19144] = 16'h3ef4;
mem_array[19147] = 16'hf433;
mem_array[19146] = 16'h3de5;
mem_array[19149] = 16'h24b5;
mem_array[19148] = 16'h3d89;
mem_array[19151] = 16'h9dbd;
mem_array[19150] = 16'h3d2d;
mem_array[19153] = 16'hef36;
mem_array[19152] = 16'h3d9f;
mem_array[19155] = 16'h387d;
mem_array[19154] = 16'h3e6b;
mem_array[19157] = 16'h1635;
mem_array[19156] = 16'h3f23;
mem_array[19159] = 16'h3047;
mem_array[19158] = 16'hbe3e;
mem_array[19161] = 16'h21c0;
mem_array[19160] = 16'h3d41;
mem_array[19163] = 16'hda30;
mem_array[19162] = 16'h3cf8;
mem_array[19165] = 16'h6300;
mem_array[19164] = 16'hbe53;
mem_array[19167] = 16'hfdd1;
mem_array[19166] = 16'hbf51;
mem_array[19169] = 16'hca4e;
mem_array[19168] = 16'h3ee5;
mem_array[19171] = 16'ha9b9;
mem_array[19170] = 16'hbd33;
mem_array[19173] = 16'h96bd;
mem_array[19172] = 16'h3e29;
mem_array[19175] = 16'hcd8d;
mem_array[19174] = 16'h3dd1;
mem_array[19177] = 16'ha4ba;
mem_array[19176] = 16'h3de2;
mem_array[19179] = 16'hd16a;
mem_array[19178] = 16'h3e20;
mem_array[19181] = 16'h954d;
mem_array[19180] = 16'hbe13;
mem_array[19183] = 16'h96d1;
mem_array[19182] = 16'hbd8f;
mem_array[19185] = 16'h25b7;
mem_array[19184] = 16'h3dac;
mem_array[19187] = 16'ha3b6;
mem_array[19186] = 16'h3d22;
mem_array[19189] = 16'h04a4;
mem_array[19188] = 16'hc02c;
mem_array[19191] = 16'hb2ca;
mem_array[19190] = 16'h3ec0;
mem_array[19193] = 16'hd3de;
mem_array[19192] = 16'h3db2;
mem_array[19195] = 16'h25f9;
mem_array[19194] = 16'hbd7b;
mem_array[19197] = 16'h79ce;
mem_array[19196] = 16'hbf3f;
mem_array[19199] = 16'hccf9;
mem_array[19198] = 16'hbd48;
mem_array[19201] = 16'h19c1;
mem_array[19200] = 16'h3e0a;
mem_array[19203] = 16'h1723;
mem_array[19202] = 16'h3ef8;
mem_array[19205] = 16'h1381;
mem_array[19204] = 16'hbf34;
mem_array[19207] = 16'hd1fd;
mem_array[19206] = 16'hbee2;
mem_array[19209] = 16'h7282;
mem_array[19208] = 16'h3e28;
mem_array[19211] = 16'h1b69;
mem_array[19210] = 16'h3e63;
mem_array[19213] = 16'h2059;
mem_array[19212] = 16'h3f0a;
mem_array[19215] = 16'h66f7;
mem_array[19214] = 16'h3dc1;
mem_array[19217] = 16'hd256;
mem_array[19216] = 16'h3eb8;
mem_array[19219] = 16'h1ec4;
mem_array[19218] = 16'hbddd;
mem_array[19221] = 16'hdecb;
mem_array[19220] = 16'hbde5;
mem_array[19223] = 16'hc0b7;
mem_array[19222] = 16'h3b04;
mem_array[19225] = 16'he530;
mem_array[19224] = 16'hbeee;
mem_array[19227] = 16'h0d79;
mem_array[19226] = 16'hbfa4;
mem_array[19229] = 16'h1677;
mem_array[19228] = 16'h3efb;
mem_array[19231] = 16'hac4f;
mem_array[19230] = 16'hbd28;
mem_array[19233] = 16'h46c6;
mem_array[19232] = 16'hbe1b;
mem_array[19235] = 16'hcbe7;
mem_array[19234] = 16'h3ea3;
mem_array[19237] = 16'he8d7;
mem_array[19236] = 16'h3b86;
mem_array[19239] = 16'h3c7c;
mem_array[19238] = 16'h3ec4;
mem_array[19241] = 16'h1d4b;
mem_array[19240] = 16'h3e5a;
mem_array[19243] = 16'hfd09;
mem_array[19242] = 16'h3e79;
mem_array[19245] = 16'h4ae1;
mem_array[19244] = 16'h3e61;
mem_array[19247] = 16'hb2d2;
mem_array[19246] = 16'h3dbc;
mem_array[19249] = 16'h2465;
mem_array[19248] = 16'hbfe2;
mem_array[19251] = 16'h27d5;
mem_array[19250] = 16'hbdda;
mem_array[19253] = 16'hd51a;
mem_array[19252] = 16'hbd27;
mem_array[19255] = 16'hdfce;
mem_array[19254] = 16'h3e23;
mem_array[19257] = 16'h42d0;
mem_array[19256] = 16'hbf20;
mem_array[19259] = 16'h7ad7;
mem_array[19258] = 16'h3e37;
mem_array[19261] = 16'hd353;
mem_array[19260] = 16'hbef4;
mem_array[19263] = 16'h39c1;
mem_array[19262] = 16'h3d16;
mem_array[19265] = 16'h6cf8;
mem_array[19264] = 16'hbfa4;
mem_array[19267] = 16'hcd02;
mem_array[19266] = 16'hbdd5;
mem_array[19269] = 16'hae8b;
mem_array[19268] = 16'h3e30;
mem_array[19271] = 16'hdeb5;
mem_array[19270] = 16'h3ea8;
mem_array[19273] = 16'hd78f;
mem_array[19272] = 16'h3e9a;
mem_array[19275] = 16'h6737;
mem_array[19274] = 16'h3e91;
mem_array[19277] = 16'h3739;
mem_array[19276] = 16'h3d9b;
mem_array[19279] = 16'heb0c;
mem_array[19278] = 16'h3ea0;
mem_array[19281] = 16'h5c3f;
mem_array[19280] = 16'hbc48;
mem_array[19283] = 16'hd721;
mem_array[19282] = 16'hbc83;
mem_array[19285] = 16'h52d7;
mem_array[19284] = 16'hbe05;
mem_array[19287] = 16'hf47b;
mem_array[19286] = 16'hbf80;
mem_array[19289] = 16'hd486;
mem_array[19288] = 16'h3c56;
mem_array[19291] = 16'ha4bc;
mem_array[19290] = 16'hbe14;
mem_array[19293] = 16'h76a8;
mem_array[19292] = 16'hbeb0;
mem_array[19295] = 16'h69ce;
mem_array[19294] = 16'hbf93;
mem_array[19297] = 16'h763f;
mem_array[19296] = 16'hbe10;
mem_array[19299] = 16'he68d;
mem_array[19298] = 16'h3e10;
mem_array[19301] = 16'h4969;
mem_array[19300] = 16'hbe88;
mem_array[19303] = 16'h483a;
mem_array[19302] = 16'h3e14;
mem_array[19305] = 16'hfe24;
mem_array[19304] = 16'hbd51;
mem_array[19307] = 16'h7765;
mem_array[19306] = 16'h3e88;
mem_array[19309] = 16'hbb91;
mem_array[19308] = 16'hbeb4;
mem_array[19311] = 16'h5e01;
mem_array[19310] = 16'hbef4;
mem_array[19313] = 16'h277b;
mem_array[19312] = 16'hbd6b;
mem_array[19315] = 16'hcc0a;
mem_array[19314] = 16'h3d4d;
mem_array[19317] = 16'h786d;
mem_array[19316] = 16'hbece;
mem_array[19319] = 16'haa6d;
mem_array[19318] = 16'hbe55;
mem_array[19321] = 16'h02ab;
mem_array[19320] = 16'h3e2d;
mem_array[19323] = 16'ha5ec;
mem_array[19322] = 16'hbd71;
mem_array[19325] = 16'h55d2;
mem_array[19324] = 16'hbf08;
mem_array[19327] = 16'h4723;
mem_array[19326] = 16'hbead;
mem_array[19329] = 16'h2e93;
mem_array[19328] = 16'hbefa;
mem_array[19331] = 16'h6a6e;
mem_array[19330] = 16'hbd9d;
mem_array[19333] = 16'h5c74;
mem_array[19332] = 16'h3ebc;
mem_array[19335] = 16'he100;
mem_array[19334] = 16'h3ec3;
mem_array[19337] = 16'h9912;
mem_array[19336] = 16'h3e77;
mem_array[19339] = 16'he83c;
mem_array[19338] = 16'h3e9e;
mem_array[19341] = 16'h301e;
mem_array[19340] = 16'h3d06;
mem_array[19343] = 16'hf55c;
mem_array[19342] = 16'hbda3;
mem_array[19345] = 16'h599c;
mem_array[19344] = 16'hbe83;
mem_array[19347] = 16'h8d54;
mem_array[19346] = 16'hbe45;
mem_array[19349] = 16'hcfb0;
mem_array[19348] = 16'hbebc;
mem_array[19351] = 16'he532;
mem_array[19350] = 16'h3e4c;
mem_array[19353] = 16'hc0a5;
mem_array[19352] = 16'hbddd;
mem_array[19355] = 16'hdedf;
mem_array[19354] = 16'hbf94;
mem_array[19357] = 16'h6760;
mem_array[19356] = 16'h3e17;
mem_array[19359] = 16'hf97a;
mem_array[19358] = 16'hbf00;
mem_array[19361] = 16'h68d9;
mem_array[19360] = 16'hbe6a;
mem_array[19363] = 16'hc963;
mem_array[19362] = 16'h3d46;
mem_array[19365] = 16'hb1b3;
mem_array[19364] = 16'hbe48;
mem_array[19367] = 16'h45b7;
mem_array[19366] = 16'h3d10;
mem_array[19369] = 16'hfc22;
mem_array[19368] = 16'hbe02;
mem_array[19371] = 16'hffeb;
mem_array[19370] = 16'hbab5;
mem_array[19373] = 16'h68d6;
mem_array[19372] = 16'hbe17;
mem_array[19375] = 16'h1209;
mem_array[19374] = 16'hbbea;
mem_array[19377] = 16'h6526;
mem_array[19376] = 16'hbd5f;
mem_array[19379] = 16'hd7d6;
mem_array[19378] = 16'hbdde;
mem_array[19381] = 16'h0a23;
mem_array[19380] = 16'h3f24;
mem_array[19383] = 16'hb435;
mem_array[19382] = 16'hbedc;
mem_array[19385] = 16'h95d2;
mem_array[19384] = 16'h3e38;
mem_array[19387] = 16'hde8e;
mem_array[19386] = 16'hbf34;
mem_array[19389] = 16'hfe3f;
mem_array[19388] = 16'hbdf9;
mem_array[19391] = 16'h0db9;
mem_array[19390] = 16'h3e19;
mem_array[19393] = 16'hf6d2;
mem_array[19392] = 16'h3e0c;
mem_array[19395] = 16'hd359;
mem_array[19394] = 16'h3f1b;
mem_array[19397] = 16'h6eec;
mem_array[19396] = 16'hbc3f;
mem_array[19399] = 16'h7233;
mem_array[19398] = 16'h3edd;
mem_array[19401] = 16'h2c35;
mem_array[19400] = 16'hbcef;
mem_array[19403] = 16'ha427;
mem_array[19402] = 16'hbceb;
mem_array[19405] = 16'h7f72;
mem_array[19404] = 16'hbf00;
mem_array[19407] = 16'h2838;
mem_array[19406] = 16'hbf17;
mem_array[19409] = 16'ha9be;
mem_array[19408] = 16'hbeca;
mem_array[19411] = 16'hb996;
mem_array[19410] = 16'h3d31;
mem_array[19413] = 16'h8a6b;
mem_array[19412] = 16'h3e39;
mem_array[19415] = 16'hfdc2;
mem_array[19414] = 16'hbdea;
mem_array[19417] = 16'hed02;
mem_array[19416] = 16'h3eb5;
mem_array[19419] = 16'h409b;
mem_array[19418] = 16'hbf29;
mem_array[19421] = 16'h5c77;
mem_array[19420] = 16'h3d07;
mem_array[19423] = 16'h7b03;
mem_array[19422] = 16'hbda9;
mem_array[19425] = 16'h11c5;
mem_array[19424] = 16'hbf11;
mem_array[19427] = 16'hae0e;
mem_array[19426] = 16'hbe99;
mem_array[19429] = 16'h2f0e;
mem_array[19428] = 16'h3e57;
mem_array[19431] = 16'hc026;
mem_array[19430] = 16'h3de9;
mem_array[19433] = 16'h6550;
mem_array[19432] = 16'hbddb;
mem_array[19435] = 16'h6b65;
mem_array[19434] = 16'hbeb6;
mem_array[19437] = 16'hb681;
mem_array[19436] = 16'hbd85;
mem_array[19439] = 16'h423c;
mem_array[19438] = 16'hbdff;
mem_array[19441] = 16'hd6aa;
mem_array[19440] = 16'h3e64;
mem_array[19443] = 16'h2ca9;
mem_array[19442] = 16'hbe53;
mem_array[19445] = 16'h9b39;
mem_array[19444] = 16'hbe65;
mem_array[19447] = 16'h2394;
mem_array[19446] = 16'hbf7f;
mem_array[19449] = 16'h584a;
mem_array[19448] = 16'hbe18;
mem_array[19451] = 16'hf782;
mem_array[19450] = 16'hbdc2;
mem_array[19453] = 16'h6dae;
mem_array[19452] = 16'hbec0;
mem_array[19455] = 16'h2b0f;
mem_array[19454] = 16'h3e6f;
mem_array[19457] = 16'h56a2;
mem_array[19456] = 16'h3d5d;
mem_array[19459] = 16'h0ee6;
mem_array[19458] = 16'h3e66;
mem_array[19461] = 16'hf4a6;
mem_array[19460] = 16'hbb52;
mem_array[19463] = 16'he9ba;
mem_array[19462] = 16'hbddf;
mem_array[19465] = 16'h0ec0;
mem_array[19464] = 16'h3e17;
mem_array[19467] = 16'h847d;
mem_array[19466] = 16'hbec5;
mem_array[19469] = 16'hb679;
mem_array[19468] = 16'hbf1e;
mem_array[19471] = 16'h80ac;
mem_array[19470] = 16'h3e83;
mem_array[19473] = 16'h6bc2;
mem_array[19472] = 16'h3e8e;
mem_array[19475] = 16'h9ca0;
mem_array[19474] = 16'h3ece;
mem_array[19477] = 16'h3df3;
mem_array[19476] = 16'h3d95;
mem_array[19479] = 16'h0e00;
mem_array[19478] = 16'h3e80;
mem_array[19481] = 16'hae6a;
mem_array[19480] = 16'hbc91;
mem_array[19483] = 16'hf1ba;
mem_array[19482] = 16'h3eae;
mem_array[19485] = 16'h1687;
mem_array[19484] = 16'hbf4b;
mem_array[19487] = 16'hb21d;
mem_array[19486] = 16'h3ea3;
mem_array[19489] = 16'h4773;
mem_array[19488] = 16'h3d9c;
mem_array[19491] = 16'h157b;
mem_array[19490] = 16'hbd46;
mem_array[19493] = 16'h9e1a;
mem_array[19492] = 16'hbd8e;
mem_array[19495] = 16'h0288;
mem_array[19494] = 16'hbf04;
mem_array[19497] = 16'h2ab4;
mem_array[19496] = 16'h3e35;
mem_array[19499] = 16'h8482;
mem_array[19498] = 16'h3e56;
mem_array[19501] = 16'h1c8b;
mem_array[19500] = 16'h3e5c;
mem_array[19503] = 16'h4e25;
mem_array[19502] = 16'h3cd4;
mem_array[19505] = 16'ha3a5;
mem_array[19504] = 16'hbddd;
mem_array[19507] = 16'hf3ba;
mem_array[19506] = 16'hbf6c;
mem_array[19509] = 16'h6c3f;
mem_array[19508] = 16'h3e95;
mem_array[19511] = 16'hbb1c;
mem_array[19510] = 16'hbe31;
mem_array[19513] = 16'h3443;
mem_array[19512] = 16'hbe05;
mem_array[19515] = 16'h2894;
mem_array[19514] = 16'h3e22;
mem_array[19517] = 16'h1000;
mem_array[19516] = 16'h3d01;
mem_array[19519] = 16'h5ed8;
mem_array[19518] = 16'hbe8f;
mem_array[19521] = 16'h980e;
mem_array[19520] = 16'hbd81;
mem_array[19523] = 16'hd876;
mem_array[19522] = 16'h3c37;
mem_array[19525] = 16'h997e;
mem_array[19524] = 16'h3d71;
mem_array[19527] = 16'h764b;
mem_array[19526] = 16'hbeb1;
mem_array[19529] = 16'h0b1c;
mem_array[19528] = 16'hbeb9;
mem_array[19531] = 16'h5859;
mem_array[19530] = 16'h3e36;
mem_array[19533] = 16'h0740;
mem_array[19532] = 16'h3e16;
mem_array[19535] = 16'h2d04;
mem_array[19534] = 16'h3df0;
mem_array[19537] = 16'h5b14;
mem_array[19536] = 16'h3eab;
mem_array[19539] = 16'hbd57;
mem_array[19538] = 16'h3e5e;
mem_array[19541] = 16'he302;
mem_array[19540] = 16'hbdba;
mem_array[19543] = 16'hd081;
mem_array[19542] = 16'h3e94;
mem_array[19545] = 16'h6a37;
mem_array[19544] = 16'hbf24;
mem_array[19547] = 16'he71d;
mem_array[19546] = 16'h3d21;
mem_array[19549] = 16'h7ba5;
mem_array[19548] = 16'h3b63;
mem_array[19551] = 16'h4279;
mem_array[19550] = 16'h3ebb;
mem_array[19553] = 16'h82b1;
mem_array[19552] = 16'hbe8c;
mem_array[19555] = 16'h92ba;
mem_array[19554] = 16'hbf04;
mem_array[19557] = 16'hc7de;
mem_array[19556] = 16'h3e3d;
mem_array[19559] = 16'h683d;
mem_array[19558] = 16'hbc4f;
mem_array[19561] = 16'h2f97;
mem_array[19560] = 16'h3e86;
mem_array[19563] = 16'h1e80;
mem_array[19562] = 16'h3e8e;
mem_array[19565] = 16'hc3f6;
mem_array[19564] = 16'hbdf8;
mem_array[19567] = 16'hb78f;
mem_array[19566] = 16'h3e20;
mem_array[19569] = 16'h40e7;
mem_array[19568] = 16'h3e67;
mem_array[19571] = 16'h50ba;
mem_array[19570] = 16'hbf68;
mem_array[19573] = 16'hd1fb;
mem_array[19572] = 16'hbcd2;
mem_array[19575] = 16'h3f3f;
mem_array[19574] = 16'h3e3b;
mem_array[19577] = 16'h2f75;
mem_array[19576] = 16'h3d30;
mem_array[19579] = 16'hd6aa;
mem_array[19578] = 16'hbed7;
mem_array[19581] = 16'hd833;
mem_array[19580] = 16'hbd49;
mem_array[19583] = 16'h9eeb;
mem_array[19582] = 16'hbddc;
mem_array[19585] = 16'h9454;
mem_array[19584] = 16'hbd7d;
mem_array[19587] = 16'hb95c;
mem_array[19586] = 16'hbe81;
mem_array[19589] = 16'h26b6;
mem_array[19588] = 16'h3e01;
mem_array[19591] = 16'hc8b3;
mem_array[19590] = 16'h3e87;
mem_array[19593] = 16'hb3e8;
mem_array[19592] = 16'h3f00;
mem_array[19595] = 16'h2f9a;
mem_array[19594] = 16'hbb22;
mem_array[19597] = 16'h92b2;
mem_array[19596] = 16'h3d48;
mem_array[19599] = 16'hb992;
mem_array[19598] = 16'h3eb3;
mem_array[19601] = 16'hd290;
mem_array[19600] = 16'hbe63;
mem_array[19603] = 16'h89fe;
mem_array[19602] = 16'h3d1b;
mem_array[19605] = 16'h1c51;
mem_array[19604] = 16'hbe63;
mem_array[19607] = 16'h3747;
mem_array[19606] = 16'hbdcb;
mem_array[19609] = 16'he7fa;
mem_array[19608] = 16'hbd13;
mem_array[19611] = 16'h5b59;
mem_array[19610] = 16'h3df0;
mem_array[19613] = 16'hb11d;
mem_array[19612] = 16'hbdd2;
mem_array[19615] = 16'hbded;
mem_array[19614] = 16'hbf11;
mem_array[19617] = 16'h8b63;
mem_array[19616] = 16'h3d91;
mem_array[19619] = 16'hd798;
mem_array[19618] = 16'hbe94;
mem_array[19621] = 16'h311a;
mem_array[19620] = 16'hbe34;
mem_array[19623] = 16'hc482;
mem_array[19622] = 16'h3f10;
mem_array[19625] = 16'had5d;
mem_array[19624] = 16'h3e3c;
mem_array[19627] = 16'hc59c;
mem_array[19626] = 16'h3ee7;
mem_array[19629] = 16'h58ee;
mem_array[19628] = 16'hbe17;
mem_array[19631] = 16'h6f98;
mem_array[19630] = 16'hc010;
mem_array[19633] = 16'hccc2;
mem_array[19632] = 16'hbde4;
mem_array[19635] = 16'h1a33;
mem_array[19634] = 16'h3e84;
mem_array[19637] = 16'h65fd;
mem_array[19636] = 16'hbe59;
mem_array[19639] = 16'h53f0;
mem_array[19638] = 16'hbed9;
mem_array[19641] = 16'h2f1e;
mem_array[19640] = 16'hbd53;
mem_array[19643] = 16'hd469;
mem_array[19642] = 16'h3a1a;
mem_array[19645] = 16'hf8e5;
mem_array[19644] = 16'h3eac;
mem_array[19647] = 16'hc65b;
mem_array[19646] = 16'hbd09;
mem_array[19649] = 16'h0a6f;
mem_array[19648] = 16'h3e4a;
mem_array[19651] = 16'h3841;
mem_array[19650] = 16'h3e43;
mem_array[19653] = 16'hb285;
mem_array[19652] = 16'hbe83;
mem_array[19655] = 16'h99ab;
mem_array[19654] = 16'hbdd1;
mem_array[19657] = 16'hcaf1;
mem_array[19656] = 16'h3da7;
mem_array[19659] = 16'he3fc;
mem_array[19658] = 16'h3dd6;
mem_array[19661] = 16'he80a;
mem_array[19660] = 16'hbe9d;
mem_array[19663] = 16'h5de2;
mem_array[19662] = 16'hbe4a;
mem_array[19665] = 16'h6c3b;
mem_array[19664] = 16'h3e34;
mem_array[19667] = 16'hddc7;
mem_array[19666] = 16'h3e59;
mem_array[19669] = 16'h0438;
mem_array[19668] = 16'hbe2a;
mem_array[19671] = 16'h5a89;
mem_array[19670] = 16'h3ea4;
mem_array[19673] = 16'hc245;
mem_array[19672] = 16'hbe67;
mem_array[19675] = 16'h9dff;
mem_array[19674] = 16'hbf06;
mem_array[19677] = 16'h1917;
mem_array[19676] = 16'h3e81;
mem_array[19679] = 16'h253b;
mem_array[19678] = 16'hbf30;
mem_array[19681] = 16'hd2e2;
mem_array[19680] = 16'h3e73;
mem_array[19683] = 16'h4367;
mem_array[19682] = 16'h3e21;
mem_array[19685] = 16'hee60;
mem_array[19684] = 16'h3dad;
mem_array[19687] = 16'hbc58;
mem_array[19686] = 16'h3d90;
mem_array[19689] = 16'h71e2;
mem_array[19688] = 16'h3e63;
mem_array[19691] = 16'h4a14;
mem_array[19690] = 16'hc00d;
mem_array[19693] = 16'hbbc6;
mem_array[19692] = 16'hbe63;
mem_array[19695] = 16'hf337;
mem_array[19694] = 16'h3e5b;
mem_array[19697] = 16'he59d;
mem_array[19696] = 16'hbedd;
mem_array[19699] = 16'hdb1e;
mem_array[19698] = 16'hbe58;
mem_array[19701] = 16'h3cb0;
mem_array[19700] = 16'hbdbe;
mem_array[19703] = 16'hd561;
mem_array[19702] = 16'hbd89;
mem_array[19705] = 16'h329c;
mem_array[19704] = 16'hbe80;
mem_array[19707] = 16'h42cd;
mem_array[19706] = 16'h3e32;
mem_array[19709] = 16'ha4a7;
mem_array[19708] = 16'h3cb2;
mem_array[19711] = 16'h12b4;
mem_array[19710] = 16'h3e38;
mem_array[19713] = 16'he1e2;
mem_array[19712] = 16'hbe56;
mem_array[19715] = 16'h20a5;
mem_array[19714] = 16'hbe69;
mem_array[19717] = 16'hee8a;
mem_array[19716] = 16'h3e0d;
mem_array[19719] = 16'h9beb;
mem_array[19718] = 16'h3db3;
mem_array[19721] = 16'h5778;
mem_array[19720] = 16'hbe6d;
mem_array[19723] = 16'h2045;
mem_array[19722] = 16'hbca5;
mem_array[19725] = 16'h2e3a;
mem_array[19724] = 16'hbede;
mem_array[19727] = 16'h35f1;
mem_array[19726] = 16'h3c81;
mem_array[19729] = 16'h32f0;
mem_array[19728] = 16'h3ebe;
mem_array[19731] = 16'h907b;
mem_array[19730] = 16'h3eb0;
mem_array[19733] = 16'h7549;
mem_array[19732] = 16'hbef8;
mem_array[19735] = 16'hcfe0;
mem_array[19734] = 16'hbe1b;
mem_array[19737] = 16'h6c68;
mem_array[19736] = 16'hbcaf;
mem_array[19739] = 16'h8ca0;
mem_array[19738] = 16'hbf27;
mem_array[19741] = 16'hbe70;
mem_array[19740] = 16'h3d5f;
mem_array[19743] = 16'hf667;
mem_array[19742] = 16'hbdef;
mem_array[19745] = 16'hca50;
mem_array[19744] = 16'hbec9;
mem_array[19747] = 16'h7f18;
mem_array[19746] = 16'h3d96;
mem_array[19749] = 16'hf526;
mem_array[19748] = 16'hbcd7;
mem_array[19751] = 16'h3bc6;
mem_array[19750] = 16'hbfdc;
mem_array[19753] = 16'h6194;
mem_array[19752] = 16'hbf0c;
mem_array[19755] = 16'h355e;
mem_array[19754] = 16'h3e3d;
mem_array[19757] = 16'hb2b3;
mem_array[19756] = 16'h3da5;
mem_array[19759] = 16'hc6ca;
mem_array[19758] = 16'h3d9d;
mem_array[19761] = 16'he099;
mem_array[19760] = 16'h3d6c;
mem_array[19763] = 16'h6db6;
mem_array[19762] = 16'hbb4d;
mem_array[19765] = 16'h1385;
mem_array[19764] = 16'h3e4e;
mem_array[19767] = 16'h3d47;
mem_array[19766] = 16'hbe52;
mem_array[19769] = 16'h34e7;
mem_array[19768] = 16'h3d3f;
mem_array[19771] = 16'h4a42;
mem_array[19770] = 16'h3ee8;
mem_array[19773] = 16'h39a7;
mem_array[19772] = 16'hbee7;
mem_array[19775] = 16'h6d95;
mem_array[19774] = 16'hbe91;
mem_array[19777] = 16'h50e1;
mem_array[19776] = 16'h3e80;
mem_array[19779] = 16'h0415;
mem_array[19778] = 16'h3e2f;
mem_array[19781] = 16'h184a;
mem_array[19780] = 16'h3e95;
mem_array[19783] = 16'hd490;
mem_array[19782] = 16'hbd54;
mem_array[19785] = 16'hf320;
mem_array[19784] = 16'hbf14;
mem_array[19787] = 16'h93ac;
mem_array[19786] = 16'h3eb3;
mem_array[19789] = 16'he58b;
mem_array[19788] = 16'h3dd3;
mem_array[19791] = 16'h2373;
mem_array[19790] = 16'hbee4;
mem_array[19793] = 16'h3ffd;
mem_array[19792] = 16'hbf0f;
mem_array[19795] = 16'he032;
mem_array[19794] = 16'h3e26;
mem_array[19797] = 16'hdb46;
mem_array[19796] = 16'hbdd1;
mem_array[19799] = 16'h69ae;
mem_array[19798] = 16'hbe96;
mem_array[19801] = 16'h3ce8;
mem_array[19800] = 16'hbf59;
mem_array[19803] = 16'hf03c;
mem_array[19802] = 16'h3e06;
mem_array[19805] = 16'h1bd1;
mem_array[19804] = 16'h3e1f;
mem_array[19807] = 16'h23f4;
mem_array[19806] = 16'h3ec4;
mem_array[19809] = 16'hff18;
mem_array[19808] = 16'hbd2d;
mem_array[19811] = 16'h8e59;
mem_array[19810] = 16'hbf93;
mem_array[19813] = 16'hb87b;
mem_array[19812] = 16'hbf90;
mem_array[19815] = 16'he801;
mem_array[19814] = 16'h3ce6;
mem_array[19817] = 16'h24d0;
mem_array[19816] = 16'hbe46;
mem_array[19819] = 16'hca94;
mem_array[19818] = 16'h3eb7;
mem_array[19821] = 16'hbfd2;
mem_array[19820] = 16'hbddb;
mem_array[19823] = 16'h0ba7;
mem_array[19822] = 16'h3d4b;
mem_array[19825] = 16'hdc7a;
mem_array[19824] = 16'h3d82;
mem_array[19827] = 16'h3305;
mem_array[19826] = 16'hbd32;
mem_array[19829] = 16'h77fb;
mem_array[19828] = 16'h3dd7;
mem_array[19831] = 16'h38d1;
mem_array[19830] = 16'h3f3e;
mem_array[19833] = 16'hff73;
mem_array[19832] = 16'hbfac;
mem_array[19835] = 16'h44eb;
mem_array[19834] = 16'hbe45;
mem_array[19837] = 16'h6e5b;
mem_array[19836] = 16'h3e5f;
mem_array[19839] = 16'hfbcd;
mem_array[19838] = 16'hbd42;
mem_array[19841] = 16'h83a5;
mem_array[19840] = 16'h3a18;
mem_array[19843] = 16'hdf48;
mem_array[19842] = 16'hbe5e;
mem_array[19845] = 16'h6293;
mem_array[19844] = 16'hbf05;
mem_array[19847] = 16'h892a;
mem_array[19846] = 16'h3e88;
mem_array[19849] = 16'h3210;
mem_array[19848] = 16'hbf14;
mem_array[19851] = 16'hd313;
mem_array[19850] = 16'hbf08;
mem_array[19853] = 16'h71b0;
mem_array[19852] = 16'hbedc;
mem_array[19855] = 16'heab6;
mem_array[19854] = 16'h3f5e;
mem_array[19857] = 16'h7ff0;
mem_array[19856] = 16'hbe8c;
mem_array[19859] = 16'h27f0;
mem_array[19858] = 16'hbf3d;
mem_array[19861] = 16'hf807;
mem_array[19860] = 16'hbed9;
mem_array[19863] = 16'h51d0;
mem_array[19862] = 16'h3ece;
mem_array[19865] = 16'h6156;
mem_array[19864] = 16'h3dec;
mem_array[19867] = 16'h6814;
mem_array[19866] = 16'h3f10;
mem_array[19869] = 16'h3671;
mem_array[19868] = 16'h3db8;
mem_array[19871] = 16'hdb23;
mem_array[19870] = 16'hbf29;
mem_array[19873] = 16'h742a;
mem_array[19872] = 16'hbf3e;
mem_array[19875] = 16'h6f58;
mem_array[19874] = 16'h3dea;
mem_array[19877] = 16'h91f6;
mem_array[19876] = 16'hbf4f;
mem_array[19879] = 16'haa89;
mem_array[19878] = 16'h3f15;
mem_array[19881] = 16'h7e30;
mem_array[19880] = 16'h3d89;
mem_array[19883] = 16'h6121;
mem_array[19882] = 16'hbca7;
mem_array[19885] = 16'hdc52;
mem_array[19884] = 16'hbdc7;
mem_array[19887] = 16'h8755;
mem_array[19886] = 16'h3e42;
mem_array[19889] = 16'h7523;
mem_array[19888] = 16'h3dbe;
mem_array[19891] = 16'he556;
mem_array[19890] = 16'h3e81;
mem_array[19893] = 16'h8cd0;
mem_array[19892] = 16'hbf0e;
mem_array[19895] = 16'h466b;
mem_array[19894] = 16'hbefc;
mem_array[19897] = 16'hfb8b;
mem_array[19896] = 16'hbe0e;
mem_array[19899] = 16'hcc87;
mem_array[19898] = 16'hbe0c;
mem_array[19901] = 16'h6bc6;
mem_array[19900] = 16'hbf4d;
mem_array[19903] = 16'h1fc5;
mem_array[19902] = 16'hbd1c;
mem_array[19905] = 16'hcf7a;
mem_array[19904] = 16'h3e00;
mem_array[19907] = 16'ha1b2;
mem_array[19906] = 16'h3e7b;
mem_array[19909] = 16'h87d7;
mem_array[19908] = 16'hbeab;
mem_array[19911] = 16'hc97b;
mem_array[19910] = 16'hbe49;
mem_array[19913] = 16'h1ccd;
mem_array[19912] = 16'h3da0;
mem_array[19915] = 16'hddec;
mem_array[19914] = 16'h3fb6;
mem_array[19917] = 16'h1b09;
mem_array[19916] = 16'hbf67;
mem_array[19919] = 16'hc610;
mem_array[19918] = 16'hbfa1;
mem_array[19921] = 16'hfd3e;
mem_array[19920] = 16'hbee8;
mem_array[19923] = 16'h7c02;
mem_array[19922] = 16'hbea8;
mem_array[19925] = 16'ha1ef;
mem_array[19924] = 16'h3da5;
mem_array[19927] = 16'hbbe0;
mem_array[19926] = 16'h3e47;
mem_array[19929] = 16'h251b;
mem_array[19928] = 16'hbe50;
mem_array[19931] = 16'h60e6;
mem_array[19930] = 16'hbe17;
mem_array[19933] = 16'hf790;
mem_array[19932] = 16'h3d90;
mem_array[19935] = 16'heac5;
mem_array[19934] = 16'h3df2;
mem_array[19937] = 16'h3569;
mem_array[19936] = 16'h3d31;
mem_array[19939] = 16'h0539;
mem_array[19938] = 16'hbe8a;
mem_array[19941] = 16'h7b1f;
mem_array[19940] = 16'hbce0;
mem_array[19943] = 16'ha556;
mem_array[19942] = 16'h3d4b;
mem_array[19945] = 16'ha37c;
mem_array[19944] = 16'hbf66;
mem_array[19947] = 16'hcc6c;
mem_array[19946] = 16'hbe3c;
mem_array[19949] = 16'h1fa5;
mem_array[19948] = 16'hbef7;
mem_array[19951] = 16'haba9;
mem_array[19950] = 16'h3f29;
mem_array[19953] = 16'h4d3f;
mem_array[19952] = 16'hbf0e;
mem_array[19955] = 16'h2bc6;
mem_array[19954] = 16'hbf40;
mem_array[19957] = 16'h42c2;
mem_array[19956] = 16'hbf4f;
mem_array[19959] = 16'h50fc;
mem_array[19958] = 16'hbf96;
mem_array[19961] = 16'h60d9;
mem_array[19960] = 16'hbf99;
mem_array[19963] = 16'h85db;
mem_array[19962] = 16'h3ed6;
mem_array[19965] = 16'h37b5;
mem_array[19964] = 16'hbf13;
mem_array[19967] = 16'h47d4;
mem_array[19966] = 16'h3ea6;
mem_array[19969] = 16'h437a;
mem_array[19968] = 16'hbee5;
mem_array[19971] = 16'h1e48;
mem_array[19970] = 16'hbeeb;
mem_array[19973] = 16'hb4ef;
mem_array[19972] = 16'h3e69;
mem_array[19975] = 16'hcf92;
mem_array[19974] = 16'h3f7a;
mem_array[19977] = 16'hbd18;
mem_array[19976] = 16'hbeff;
mem_array[19979] = 16'hab38;
mem_array[19978] = 16'hbf9c;
mem_array[19981] = 16'h46fc;
mem_array[19980] = 16'h3eaa;
mem_array[19983] = 16'h774c;
mem_array[19982] = 16'hbeed;
mem_array[19985] = 16'hf600;
mem_array[19984] = 16'hbddc;
mem_array[19987] = 16'h14d0;
mem_array[19986] = 16'hbf66;
mem_array[19989] = 16'h2e5c;
mem_array[19988] = 16'hbf24;
mem_array[19991] = 16'h1410;
mem_array[19990] = 16'hbf18;
mem_array[19993] = 16'h77b2;
mem_array[19992] = 16'h3eba;
mem_array[19995] = 16'h5760;
mem_array[19994] = 16'h3f1c;
mem_array[19997] = 16'h78c6;
mem_array[19996] = 16'h3f62;
mem_array[19999] = 16'h997b;
mem_array[19998] = 16'h3d54;
mem_array[20001] = 16'h00c0;
mem_array[20000] = 16'h3d6b;
mem_array[20003] = 16'h578b;
mem_array[20002] = 16'hbd0d;
mem_array[20005] = 16'hd86f;
mem_array[20004] = 16'hbf71;
mem_array[20007] = 16'h7c53;
mem_array[20006] = 16'hbe98;
mem_array[20009] = 16'hb245;
mem_array[20008] = 16'h3d4c;
mem_array[20011] = 16'h80ac;
mem_array[20010] = 16'hbe90;
mem_array[20013] = 16'h1b69;
mem_array[20012] = 16'h3f38;
mem_array[20015] = 16'h9a28;
mem_array[20014] = 16'hbe38;
mem_array[20017] = 16'h8f25;
mem_array[20016] = 16'hbeeb;
mem_array[20019] = 16'h090a;
mem_array[20018] = 16'hbf19;
mem_array[20021] = 16'hd1e7;
mem_array[20020] = 16'hbf61;
mem_array[20023] = 16'h5886;
mem_array[20022] = 16'h3f48;
mem_array[20025] = 16'h6230;
mem_array[20024] = 16'hbf44;
mem_array[20027] = 16'h5ffc;
mem_array[20026] = 16'hbe9f;
mem_array[20029] = 16'ha5a1;
mem_array[20028] = 16'hbf30;
mem_array[20031] = 16'h7ec6;
mem_array[20030] = 16'hbebd;
mem_array[20033] = 16'h1f0d;
mem_array[20032] = 16'h3f1b;
mem_array[20035] = 16'h0c43;
mem_array[20034] = 16'h4008;
mem_array[20037] = 16'hfd43;
mem_array[20036] = 16'h3ca5;
mem_array[20039] = 16'h5520;
mem_array[20038] = 16'hbf3b;
mem_array[20041] = 16'h0624;
mem_array[20040] = 16'h3eb0;
mem_array[20043] = 16'h26ee;
mem_array[20042] = 16'hbf26;
mem_array[20045] = 16'hd89a;
mem_array[20044] = 16'hbf87;
mem_array[20047] = 16'h7e55;
mem_array[20046] = 16'hbfc6;
mem_array[20049] = 16'hddf1;
mem_array[20048] = 16'hbf57;
mem_array[20051] = 16'h3c6c;
mem_array[20050] = 16'h3eed;
mem_array[20053] = 16'h7c7a;
mem_array[20052] = 16'hbf02;
mem_array[20055] = 16'h1fa0;
mem_array[20054] = 16'hbfac;
mem_array[20057] = 16'haf30;
mem_array[20056] = 16'hbf77;
mem_array[20059] = 16'h14ee;
mem_array[20058] = 16'h3eb2;
mem_array[20061] = 16'h920c;
mem_array[20060] = 16'h3c87;
mem_array[20063] = 16'h3348;
mem_array[20062] = 16'hbcd4;
mem_array[20065] = 16'hd58b;
mem_array[20064] = 16'hbf79;
mem_array[20067] = 16'h5724;
mem_array[20066] = 16'hbfe3;
mem_array[20069] = 16'h8f83;
mem_array[20068] = 16'h3e70;
mem_array[20071] = 16'h3048;
mem_array[20070] = 16'h3fb1;
mem_array[20073] = 16'h9ff0;
mem_array[20072] = 16'hbedc;
mem_array[20075] = 16'h2c16;
mem_array[20074] = 16'hbd90;
mem_array[20077] = 16'h0e7c;
mem_array[20076] = 16'hbf95;
mem_array[20079] = 16'h3fab;
mem_array[20078] = 16'h3e81;
mem_array[20081] = 16'h8143;
mem_array[20080] = 16'hbfee;
mem_array[20083] = 16'hca80;
mem_array[20082] = 16'hbeda;
mem_array[20085] = 16'h1ea0;
mem_array[20084] = 16'h3e30;
mem_array[20087] = 16'hd9fe;
mem_array[20086] = 16'hbf89;
mem_array[20089] = 16'hebcd;
mem_array[20088] = 16'hbf61;
mem_array[20091] = 16'h1515;
mem_array[20090] = 16'hbf0a;
mem_array[20093] = 16'hd294;
mem_array[20092] = 16'h3fa4;
mem_array[20095] = 16'haa3f;
mem_array[20094] = 16'h3f75;
mem_array[20097] = 16'h66da;
mem_array[20096] = 16'h3f10;
mem_array[20099] = 16'h9afe;
mem_array[20098] = 16'hbf32;
mem_array[20101] = 16'h5da6;
mem_array[20100] = 16'h3ed3;
mem_array[20103] = 16'h6cb0;
mem_array[20102] = 16'hbe6f;
mem_array[20105] = 16'h6ce9;
mem_array[20104] = 16'hbe4c;
mem_array[20107] = 16'h57e7;
mem_array[20106] = 16'h3def;
mem_array[20109] = 16'h57d0;
mem_array[20108] = 16'h3e18;
mem_array[20111] = 16'h7cce;
mem_array[20110] = 16'h3f03;
mem_array[20113] = 16'h048c;
mem_array[20112] = 16'hbe95;
mem_array[20115] = 16'h5033;
mem_array[20114] = 16'hbce1;
mem_array[20117] = 16'h6e08;
mem_array[20116] = 16'h3e13;
mem_array[20119] = 16'hf9d8;
mem_array[20118] = 16'h3f89;
mem_array[20121] = 16'h5ca7;
mem_array[20120] = 16'h3dd1;
mem_array[20123] = 16'ha64d;
mem_array[20122] = 16'hbd99;
mem_array[20125] = 16'h704f;
mem_array[20124] = 16'hbdc1;
mem_array[20127] = 16'h60d2;
mem_array[20126] = 16'hbddf;
mem_array[20129] = 16'hbf36;
mem_array[20128] = 16'hbd28;
mem_array[20131] = 16'h25f1;
mem_array[20130] = 16'hbd79;
mem_array[20133] = 16'h534b;
mem_array[20132] = 16'hbd89;
mem_array[20135] = 16'h4fa6;
mem_array[20134] = 16'hbe04;
mem_array[20137] = 16'h874b;
mem_array[20136] = 16'hbd18;
mem_array[20139] = 16'h9527;
mem_array[20138] = 16'h3e59;
mem_array[20141] = 16'h172e;
mem_array[20140] = 16'h3a1b;
mem_array[20143] = 16'h6d91;
mem_array[20142] = 16'hbe44;
mem_array[20145] = 16'hef3a;
mem_array[20144] = 16'h3bb3;
mem_array[20147] = 16'h1454;
mem_array[20146] = 16'hbeff;
mem_array[20149] = 16'h7eea;
mem_array[20148] = 16'hbeed;
mem_array[20151] = 16'h46d1;
mem_array[20150] = 16'h3c32;
mem_array[20153] = 16'h500e;
mem_array[20152] = 16'hbe48;
mem_array[20155] = 16'h4044;
mem_array[20154] = 16'hbe67;
mem_array[20157] = 16'h9bbd;
mem_array[20156] = 16'h3cbf;
mem_array[20159] = 16'h1f4a;
mem_array[20158] = 16'h3cfb;
mem_array[20161] = 16'he988;
mem_array[20160] = 16'hbd49;
mem_array[20163] = 16'h387a;
mem_array[20162] = 16'hbd8b;
mem_array[20165] = 16'h0428;
mem_array[20164] = 16'hbd03;
mem_array[20167] = 16'h7032;
mem_array[20166] = 16'h3c4c;
mem_array[20169] = 16'h5208;
mem_array[20168] = 16'h3cd2;
mem_array[20171] = 16'hd7af;
mem_array[20170] = 16'h3d24;
mem_array[20173] = 16'hc1a7;
mem_array[20172] = 16'hbd14;
mem_array[20175] = 16'h8294;
mem_array[20174] = 16'hbd29;
mem_array[20177] = 16'ha641;
mem_array[20176] = 16'h3caa;
mem_array[20179] = 16'h5c85;
mem_array[20178] = 16'hbd2e;
mem_array[20181] = 16'h75f9;
mem_array[20180] = 16'hbd4d;
mem_array[20183] = 16'hf511;
mem_array[20182] = 16'h3d81;
mem_array[20185] = 16'hde04;
mem_array[20184] = 16'hbdb7;
mem_array[20187] = 16'h20e1;
mem_array[20186] = 16'hbc77;
mem_array[20189] = 16'hb544;
mem_array[20188] = 16'hbc50;
mem_array[20191] = 16'h8303;
mem_array[20190] = 16'h3d09;
mem_array[20193] = 16'haf0b;
mem_array[20192] = 16'h3de4;
mem_array[20195] = 16'hdcb8;
mem_array[20194] = 16'h3bfd;
mem_array[20197] = 16'h1447;
mem_array[20196] = 16'h3cd9;
mem_array[20199] = 16'h7f15;
mem_array[20198] = 16'h3dbc;
mem_array[20201] = 16'h5bcb;
mem_array[20200] = 16'hbe03;
mem_array[20203] = 16'h6005;
mem_array[20202] = 16'h3d32;
mem_array[20205] = 16'h4e69;
mem_array[20204] = 16'hbd98;
mem_array[20207] = 16'hec44;
mem_array[20206] = 16'hbb74;
mem_array[20209] = 16'h5299;
mem_array[20208] = 16'hbccd;
mem_array[20211] = 16'h4b68;
mem_array[20210] = 16'h3c5e;
mem_array[20213] = 16'h10bc;
mem_array[20212] = 16'hbdba;
mem_array[20215] = 16'h0de7;
mem_array[20214] = 16'h3d63;
mem_array[20217] = 16'h1a0f;
mem_array[20216] = 16'hbd93;
mem_array[20219] = 16'h7c3e;
mem_array[20218] = 16'hbcc4;
mem_array[20221] = 16'h21bd;
mem_array[20220] = 16'hbcd8;
mem_array[20223] = 16'h5572;
mem_array[20222] = 16'h3ec9;
mem_array[20225] = 16'hac3d;
mem_array[20224] = 16'h3e7c;
mem_array[20227] = 16'h64d4;
mem_array[20226] = 16'h3e5c;
mem_array[20229] = 16'h5ce9;
mem_array[20228] = 16'h3e59;
mem_array[20231] = 16'h70fc;
mem_array[20230] = 16'hbda8;
mem_array[20233] = 16'h8cfa;
mem_array[20232] = 16'h3c3b;
mem_array[20235] = 16'h148c;
mem_array[20234] = 16'h3e60;
mem_array[20237] = 16'hc4f8;
mem_array[20236] = 16'hbead;
mem_array[20239] = 16'h8cc0;
mem_array[20238] = 16'h3ea9;
mem_array[20241] = 16'hff54;
mem_array[20240] = 16'hbd31;
mem_array[20243] = 16'h1644;
mem_array[20242] = 16'h3c14;
mem_array[20245] = 16'he188;
mem_array[20244] = 16'h3f1b;
mem_array[20247] = 16'hfee2;
mem_array[20246] = 16'hbf1f;
mem_array[20249] = 16'hcdc9;
mem_array[20248] = 16'hbe16;
mem_array[20251] = 16'h7e6e;
mem_array[20250] = 16'hbe83;
mem_array[20253] = 16'h6650;
mem_array[20252] = 16'hbdf9;
mem_array[20255] = 16'hbc3e;
mem_array[20254] = 16'h3e74;
mem_array[20257] = 16'h1944;
mem_array[20256] = 16'h3f82;
mem_array[20259] = 16'h5e4f;
mem_array[20258] = 16'h3f02;
mem_array[20261] = 16'hbdbb;
mem_array[20260] = 16'hbd5c;
mem_array[20263] = 16'h06d2;
mem_array[20262] = 16'hbe69;
mem_array[20265] = 16'h9f9b;
mem_array[20264] = 16'h3da9;
mem_array[20267] = 16'hf58c;
mem_array[20266] = 16'hbf2e;
mem_array[20269] = 16'h0d63;
mem_array[20268] = 16'hbf3b;
mem_array[20271] = 16'hd7b4;
mem_array[20270] = 16'h3f6d;
mem_array[20273] = 16'h5352;
mem_array[20272] = 16'hbf18;
mem_array[20275] = 16'hea2e;
mem_array[20274] = 16'h3ec2;
mem_array[20277] = 16'h975f;
mem_array[20276] = 16'hbf23;
mem_array[20279] = 16'he873;
mem_array[20278] = 16'hbeef;
mem_array[20281] = 16'ha5cd;
mem_array[20280] = 16'hbdc6;
mem_array[20283] = 16'hcbde;
mem_array[20282] = 16'h3dfd;
mem_array[20285] = 16'h83dd;
mem_array[20284] = 16'hbd32;
mem_array[20287] = 16'hb765;
mem_array[20286] = 16'h3d7e;
mem_array[20289] = 16'heec3;
mem_array[20288] = 16'h3d93;
mem_array[20291] = 16'h90ab;
mem_array[20290] = 16'h3e86;
mem_array[20293] = 16'hcc9a;
mem_array[20292] = 16'h3da3;
mem_array[20295] = 16'h3c5a;
mem_array[20294] = 16'h3e76;
mem_array[20297] = 16'h68de;
mem_array[20296] = 16'h3e47;
mem_array[20299] = 16'h52d1;
mem_array[20298] = 16'h3f14;
mem_array[20301] = 16'h4fb8;
mem_array[20300] = 16'hbd82;
mem_array[20303] = 16'hf2d2;
mem_array[20302] = 16'h3cc7;
mem_array[20305] = 16'hf10e;
mem_array[20304] = 16'h3dd2;
mem_array[20307] = 16'he082;
mem_array[20306] = 16'hbf11;
mem_array[20309] = 16'h3327;
mem_array[20308] = 16'hbf42;
mem_array[20311] = 16'h1ed6;
mem_array[20310] = 16'h3de3;
mem_array[20313] = 16'h3806;
mem_array[20312] = 16'hbdf3;
mem_array[20315] = 16'hfba7;
mem_array[20314] = 16'hbe72;
mem_array[20317] = 16'h0310;
mem_array[20316] = 16'h3e92;
mem_array[20319] = 16'h9ed1;
mem_array[20318] = 16'hbe22;
mem_array[20321] = 16'h6419;
mem_array[20320] = 16'hbf02;
mem_array[20323] = 16'haa47;
mem_array[20322] = 16'hbe54;
mem_array[20325] = 16'h49e1;
mem_array[20324] = 16'h3d99;
mem_array[20327] = 16'hb5dc;
mem_array[20326] = 16'h3e78;
mem_array[20329] = 16'h9abb;
mem_array[20328] = 16'hbf9b;
mem_array[20331] = 16'hcedd;
mem_array[20330] = 16'h3ef5;
mem_array[20333] = 16'h0860;
mem_array[20332] = 16'hbe9d;
mem_array[20335] = 16'hbf17;
mem_array[20334] = 16'h3ed3;
mem_array[20337] = 16'h4488;
mem_array[20336] = 16'hbf02;
mem_array[20339] = 16'hf6dd;
mem_array[20338] = 16'hbec4;
mem_array[20341] = 16'hcf94;
mem_array[20340] = 16'hbbd2;
mem_array[20343] = 16'h732f;
mem_array[20342] = 16'h3f45;
mem_array[20345] = 16'ha605;
mem_array[20344] = 16'h3ec7;
mem_array[20347] = 16'h2f59;
mem_array[20346] = 16'hbf42;
mem_array[20349] = 16'h40fa;
mem_array[20348] = 16'hbe4b;
mem_array[20351] = 16'hf3a2;
mem_array[20350] = 16'h3f01;
mem_array[20353] = 16'ha801;
mem_array[20352] = 16'hbf84;
mem_array[20355] = 16'h12e6;
mem_array[20354] = 16'hbd18;
mem_array[20357] = 16'h7e4a;
mem_array[20356] = 16'h3e34;
mem_array[20359] = 16'h2e52;
mem_array[20358] = 16'hbf14;
mem_array[20361] = 16'h1b6d;
mem_array[20360] = 16'h3d1c;
mem_array[20363] = 16'h0d59;
mem_array[20362] = 16'h3cc4;
mem_array[20365] = 16'hbfcf;
mem_array[20364] = 16'hbfb1;
mem_array[20367] = 16'h812f;
mem_array[20366] = 16'hbf71;
mem_array[20369] = 16'h1838;
mem_array[20368] = 16'hbf2e;
mem_array[20371] = 16'he310;
mem_array[20370] = 16'h3da0;
mem_array[20373] = 16'h9010;
mem_array[20372] = 16'h3e09;
mem_array[20375] = 16'h621d;
mem_array[20374] = 16'h3e38;
mem_array[20377] = 16'h346e;
mem_array[20376] = 16'h3edb;
mem_array[20379] = 16'h5087;
mem_array[20378] = 16'h3ea5;
mem_array[20381] = 16'he91c;
mem_array[20380] = 16'hbf3c;
mem_array[20383] = 16'headb;
mem_array[20382] = 16'hbedd;
mem_array[20385] = 16'h1395;
mem_array[20384] = 16'hbe7a;
mem_array[20387] = 16'hf1d7;
mem_array[20386] = 16'h3c8f;
mem_array[20389] = 16'h2389;
mem_array[20388] = 16'hbe20;
mem_array[20391] = 16'hd5e2;
mem_array[20390] = 16'h3e47;
mem_array[20393] = 16'h4b36;
mem_array[20392] = 16'hbeef;
mem_array[20395] = 16'h0e63;
mem_array[20394] = 16'h3e1b;
mem_array[20397] = 16'h087a;
mem_array[20396] = 16'hbdf6;
mem_array[20399] = 16'h68b1;
mem_array[20398] = 16'h3f06;
mem_array[20401] = 16'h7113;
mem_array[20400] = 16'h3e80;
mem_array[20403] = 16'hf6cf;
mem_array[20402] = 16'hbd42;
mem_array[20405] = 16'hd820;
mem_array[20404] = 16'h3f19;
mem_array[20407] = 16'h1845;
mem_array[20406] = 16'hbe18;
mem_array[20409] = 16'h8b9b;
mem_array[20408] = 16'hbf02;
mem_array[20411] = 16'h73f9;
mem_array[20410] = 16'h3dd8;
mem_array[20413] = 16'h2a93;
mem_array[20412] = 16'hbf37;
mem_array[20415] = 16'h2b14;
mem_array[20414] = 16'h3d22;
mem_array[20417] = 16'hc9a7;
mem_array[20416] = 16'hbec8;
mem_array[20419] = 16'h37ee;
mem_array[20418] = 16'hbe20;
mem_array[20421] = 16'h6664;
mem_array[20420] = 16'hbd8d;
mem_array[20423] = 16'h8dc5;
mem_array[20422] = 16'hbd53;
mem_array[20425] = 16'h5e27;
mem_array[20424] = 16'hbf2d;
mem_array[20427] = 16'h9123;
mem_array[20426] = 16'hbfd6;
mem_array[20429] = 16'hdcb4;
mem_array[20428] = 16'hbf0b;
mem_array[20431] = 16'h45a1;
mem_array[20430] = 16'h3e29;
mem_array[20433] = 16'h04bf;
mem_array[20432] = 16'h3f58;
mem_array[20435] = 16'h27d1;
mem_array[20434] = 16'hbebc;
mem_array[20437] = 16'h2c6a;
mem_array[20436] = 16'h3e83;
mem_array[20439] = 16'h0bef;
mem_array[20438] = 16'hbee4;
mem_array[20441] = 16'h7654;
mem_array[20440] = 16'hbf71;
mem_array[20443] = 16'h5729;
mem_array[20442] = 16'h3e93;
mem_array[20445] = 16'h12d4;
mem_array[20444] = 16'hbe9b;
mem_array[20447] = 16'h4169;
mem_array[20446] = 16'h3e94;
mem_array[20449] = 16'h2631;
mem_array[20448] = 16'h3cef;
mem_array[20451] = 16'h060d;
mem_array[20450] = 16'hbea6;
mem_array[20453] = 16'h0609;
mem_array[20452] = 16'h3ea7;
mem_array[20455] = 16'hb722;
mem_array[20454] = 16'hbf97;
mem_array[20457] = 16'h7988;
mem_array[20456] = 16'hbf71;
mem_array[20459] = 16'hf5d8;
mem_array[20458] = 16'hbef9;
mem_array[20461] = 16'hbbce;
mem_array[20460] = 16'hbf14;
mem_array[20463] = 16'he573;
mem_array[20462] = 16'h3e09;
mem_array[20465] = 16'hc041;
mem_array[20464] = 16'h3ed1;
mem_array[20467] = 16'hf531;
mem_array[20466] = 16'hbeea;
mem_array[20469] = 16'h1565;
mem_array[20468] = 16'h3c7f;
mem_array[20471] = 16'h76e2;
mem_array[20470] = 16'h3e74;
mem_array[20473] = 16'h0a9f;
mem_array[20472] = 16'hbe81;
mem_array[20475] = 16'hc7ee;
mem_array[20474] = 16'h3dba;
mem_array[20477] = 16'h8c01;
mem_array[20476] = 16'h3f00;
mem_array[20479] = 16'hd9ee;
mem_array[20478] = 16'h3ed8;
mem_array[20481] = 16'h67a4;
mem_array[20480] = 16'hbdd9;
mem_array[20483] = 16'h45ba;
mem_array[20482] = 16'h3cf1;
mem_array[20485] = 16'h01dd;
mem_array[20484] = 16'hbecc;
mem_array[20487] = 16'h5695;
mem_array[20486] = 16'hbff6;
mem_array[20489] = 16'h7241;
mem_array[20488] = 16'hbf3f;
mem_array[20491] = 16'h0a31;
mem_array[20490] = 16'h3e00;
mem_array[20493] = 16'h4d94;
mem_array[20492] = 16'h3f36;
mem_array[20495] = 16'h8fb3;
mem_array[20494] = 16'h3e77;
mem_array[20497] = 16'ha6c9;
mem_array[20496] = 16'h3e81;
mem_array[20499] = 16'h3aec;
mem_array[20498] = 16'hbcac;
mem_array[20501] = 16'h9428;
mem_array[20500] = 16'hbf62;
mem_array[20503] = 16'h82a2;
mem_array[20502] = 16'hbde6;
mem_array[20505] = 16'hbb52;
mem_array[20504] = 16'hbf05;
mem_array[20507] = 16'h9cad;
mem_array[20506] = 16'hbd8c;
mem_array[20509] = 16'h2e4e;
mem_array[20508] = 16'h3e56;
mem_array[20511] = 16'h6275;
mem_array[20510] = 16'h3eac;
mem_array[20513] = 16'h4a5f;
mem_array[20512] = 16'h3d3e;
mem_array[20515] = 16'h84d2;
mem_array[20514] = 16'hbf22;
mem_array[20517] = 16'he1e6;
mem_array[20516] = 16'hbfc6;
mem_array[20519] = 16'h1b0e;
mem_array[20518] = 16'h3e3b;
mem_array[20521] = 16'h0b38;
mem_array[20520] = 16'hbe22;
mem_array[20523] = 16'h0115;
mem_array[20522] = 16'h3e28;
mem_array[20525] = 16'h139f;
mem_array[20524] = 16'h3e25;
mem_array[20527] = 16'ha936;
mem_array[20526] = 16'h3ea8;
mem_array[20529] = 16'hb501;
mem_array[20528] = 16'hbdf9;
mem_array[20531] = 16'ha1f2;
mem_array[20530] = 16'hbe33;
mem_array[20533] = 16'h9e49;
mem_array[20532] = 16'hbf61;
mem_array[20535] = 16'hb8c9;
mem_array[20534] = 16'hbe5a;
mem_array[20537] = 16'h0f9e;
mem_array[20536] = 16'hbdff;
mem_array[20539] = 16'hb98b;
mem_array[20538] = 16'hbe86;
mem_array[20541] = 16'h57cc;
mem_array[20540] = 16'hbd3f;
mem_array[20543] = 16'h827c;
mem_array[20542] = 16'hbd89;
mem_array[20545] = 16'hd16e;
mem_array[20544] = 16'hbea7;
mem_array[20547] = 16'hc34b;
mem_array[20546] = 16'hc00a;
mem_array[20549] = 16'hf54d;
mem_array[20548] = 16'hbf1d;
mem_array[20551] = 16'h71df;
mem_array[20550] = 16'hbdaf;
mem_array[20553] = 16'hbdd2;
mem_array[20552] = 16'hbef0;
mem_array[20555] = 16'h82aa;
mem_array[20554] = 16'h3e45;
mem_array[20557] = 16'h205a;
mem_array[20556] = 16'h3e08;
mem_array[20559] = 16'h7a3d;
mem_array[20558] = 16'hbe59;
mem_array[20561] = 16'h774a;
mem_array[20560] = 16'hbe0d;
mem_array[20563] = 16'h8c68;
mem_array[20562] = 16'hbcc6;
mem_array[20565] = 16'h018c;
mem_array[20564] = 16'hbd83;
mem_array[20567] = 16'h3930;
mem_array[20566] = 16'h3d8f;
mem_array[20569] = 16'he075;
mem_array[20568] = 16'hbfb4;
mem_array[20571] = 16'hd52c;
mem_array[20570] = 16'hbf0c;
mem_array[20573] = 16'he893;
mem_array[20572] = 16'hbd14;
mem_array[20575] = 16'h7b0d;
mem_array[20574] = 16'h3d9a;
mem_array[20577] = 16'h1de5;
mem_array[20576] = 16'hbfc3;
mem_array[20579] = 16'h1f94;
mem_array[20578] = 16'h3d40;
mem_array[20581] = 16'hd036;
mem_array[20580] = 16'hbf72;
mem_array[20583] = 16'hdf1f;
mem_array[20582] = 16'h3e39;
mem_array[20585] = 16'h4043;
mem_array[20584] = 16'h3d36;
mem_array[20587] = 16'hd5c6;
mem_array[20586] = 16'hbd08;
mem_array[20589] = 16'h3c44;
mem_array[20588] = 16'hbde6;
mem_array[20591] = 16'h8abd;
mem_array[20590] = 16'h3eb2;
mem_array[20593] = 16'h5144;
mem_array[20592] = 16'hbf64;
mem_array[20595] = 16'hc289;
mem_array[20594] = 16'h3ed6;
mem_array[20597] = 16'h9b4b;
mem_array[20596] = 16'hbe0d;
mem_array[20599] = 16'hb4e9;
mem_array[20598] = 16'h3d0b;
mem_array[20601] = 16'h270b;
mem_array[20600] = 16'h3d17;
mem_array[20603] = 16'h75df;
mem_array[20602] = 16'h3c6f;
mem_array[20605] = 16'hbdc0;
mem_array[20604] = 16'hbe66;
mem_array[20607] = 16'h445e;
mem_array[20606] = 16'hc007;
mem_array[20609] = 16'h3e13;
mem_array[20608] = 16'hbf7b;
mem_array[20611] = 16'h8c11;
mem_array[20610] = 16'h3d9c;
mem_array[20613] = 16'h42b5;
mem_array[20612] = 16'hbf54;
mem_array[20615] = 16'h3c86;
mem_array[20614] = 16'h3b1a;
mem_array[20617] = 16'h8578;
mem_array[20616] = 16'h3d26;
mem_array[20619] = 16'heecf;
mem_array[20618] = 16'hbdcf;
mem_array[20621] = 16'h7b6e;
mem_array[20620] = 16'h3d4f;
mem_array[20623] = 16'h0b0c;
mem_array[20622] = 16'h3d2c;
mem_array[20625] = 16'hb725;
mem_array[20624] = 16'hbf0b;
mem_array[20627] = 16'h62ec;
mem_array[20626] = 16'hbe33;
mem_array[20629] = 16'h64ca;
mem_array[20628] = 16'hc005;
mem_array[20631] = 16'h1aa9;
mem_array[20630] = 16'h3e26;
mem_array[20633] = 16'h2abb;
mem_array[20632] = 16'hbdbe;
mem_array[20635] = 16'h29a4;
mem_array[20634] = 16'hbdb6;
mem_array[20637] = 16'h1065;
mem_array[20636] = 16'hbf13;
mem_array[20639] = 16'h6519;
mem_array[20638] = 16'h3d37;
mem_array[20641] = 16'h19e1;
mem_array[20640] = 16'hbf89;
mem_array[20643] = 16'h2221;
mem_array[20642] = 16'h3dbd;
mem_array[20645] = 16'h15bf;
mem_array[20644] = 16'h3f0b;
mem_array[20647] = 16'h2b2a;
mem_array[20646] = 16'hbecb;
mem_array[20649] = 16'h027b;
mem_array[20648] = 16'hbd85;
mem_array[20651] = 16'hed44;
mem_array[20650] = 16'hbe2a;
mem_array[20653] = 16'he638;
mem_array[20652] = 16'h3dc4;
mem_array[20655] = 16'hf3d9;
mem_array[20654] = 16'h3ef1;
mem_array[20657] = 16'hefa1;
mem_array[20656] = 16'h3d33;
mem_array[20659] = 16'h413e;
mem_array[20658] = 16'h3d5c;
mem_array[20661] = 16'hb4a4;
mem_array[20660] = 16'hbcef;
mem_array[20663] = 16'hddbc;
mem_array[20662] = 16'h3c35;
mem_array[20665] = 16'hc1b0;
mem_array[20664] = 16'hbd6b;
mem_array[20667] = 16'hd59c;
mem_array[20666] = 16'hc000;
mem_array[20669] = 16'ha31c;
mem_array[20668] = 16'hbcab;
mem_array[20671] = 16'hd861;
mem_array[20670] = 16'h3e04;
mem_array[20673] = 16'hbccc;
mem_array[20672] = 16'hbf8a;
mem_array[20675] = 16'heac9;
mem_array[20674] = 16'hbe08;
mem_array[20677] = 16'h975f;
mem_array[20676] = 16'hbddc;
mem_array[20679] = 16'hc6d0;
mem_array[20678] = 16'h3e80;
mem_array[20681] = 16'h8231;
mem_array[20680] = 16'h3e23;
mem_array[20683] = 16'h3eb9;
mem_array[20682] = 16'h3e1a;
mem_array[20685] = 16'hd944;
mem_array[20684] = 16'hbc42;
mem_array[20687] = 16'hfe55;
mem_array[20686] = 16'h3d7b;
mem_array[20689] = 16'h8a6f;
mem_array[20688] = 16'hc060;
mem_array[20691] = 16'he9ed;
mem_array[20690] = 16'hbd6d;
mem_array[20693] = 16'h4fb5;
mem_array[20692] = 16'hbe16;
mem_array[20695] = 16'h7aad;
mem_array[20694] = 16'h3dfd;
mem_array[20697] = 16'ha761;
mem_array[20696] = 16'hbef8;
mem_array[20699] = 16'h420e;
mem_array[20698] = 16'h3ee5;
mem_array[20701] = 16'h96b0;
mem_array[20700] = 16'h3d84;
mem_array[20703] = 16'h3d59;
mem_array[20702] = 16'h3dad;
mem_array[20705] = 16'h4db3;
mem_array[20704] = 16'h3dca;
mem_array[20707] = 16'h9059;
mem_array[20706] = 16'hbd8e;
mem_array[20709] = 16'h04d2;
mem_array[20708] = 16'hbdb3;
mem_array[20711] = 16'h4666;
mem_array[20710] = 16'hbd65;
mem_array[20713] = 16'h2917;
mem_array[20712] = 16'h3f00;
mem_array[20715] = 16'h934c;
mem_array[20714] = 16'h3e3b;
mem_array[20717] = 16'h5940;
mem_array[20716] = 16'hbdbc;
mem_array[20719] = 16'hd415;
mem_array[20718] = 16'h3dd9;
mem_array[20721] = 16'hfdd6;
mem_array[20720] = 16'h3d21;
mem_array[20723] = 16'hc207;
mem_array[20722] = 16'hbdf1;
mem_array[20725] = 16'h950e;
mem_array[20724] = 16'hbe29;
mem_array[20727] = 16'hd973;
mem_array[20726] = 16'hc006;
mem_array[20729] = 16'hcddf;
mem_array[20728] = 16'hbe17;
mem_array[20731] = 16'hc2b9;
mem_array[20730] = 16'hbddf;
mem_array[20733] = 16'h49f3;
mem_array[20732] = 16'h3d12;
mem_array[20735] = 16'hd684;
mem_array[20734] = 16'hbd2c;
mem_array[20737] = 16'h037b;
mem_array[20736] = 16'hbdde;
mem_array[20739] = 16'hb3fd;
mem_array[20738] = 16'h3e89;
mem_array[20741] = 16'heaf3;
mem_array[20740] = 16'h3d2a;
mem_array[20743] = 16'he10f;
mem_array[20742] = 16'h3e5e;
mem_array[20745] = 16'ha458;
mem_array[20744] = 16'hbe2e;
mem_array[20747] = 16'h3e01;
mem_array[20746] = 16'h3e29;
mem_array[20749] = 16'hf63e;
mem_array[20748] = 16'hc044;
mem_array[20751] = 16'h4e28;
mem_array[20750] = 16'hbece;
mem_array[20753] = 16'h1e96;
mem_array[20752] = 16'hbcd1;
mem_array[20755] = 16'hf9e1;
mem_array[20754] = 16'h3d88;
mem_array[20757] = 16'hfc0b;
mem_array[20756] = 16'hbe69;
mem_array[20759] = 16'hc48a;
mem_array[20758] = 16'h3e4b;
mem_array[20761] = 16'hb6ed;
mem_array[20760] = 16'hbe15;
mem_array[20763] = 16'h54fe;
mem_array[20762] = 16'h3ddf;
mem_array[20765] = 16'h2bbc;
mem_array[20764] = 16'h3d2a;
mem_array[20767] = 16'h73cb;
mem_array[20766] = 16'h3d82;
mem_array[20769] = 16'h71f4;
mem_array[20768] = 16'h3d6d;
mem_array[20771] = 16'h388b;
mem_array[20770] = 16'h3e07;
mem_array[20773] = 16'h4ff7;
mem_array[20772] = 16'h3f2b;
mem_array[20775] = 16'hf5c6;
mem_array[20774] = 16'hbcf2;
mem_array[20777] = 16'h4849;
mem_array[20776] = 16'hbf1f;
mem_array[20779] = 16'hc8ec;
mem_array[20778] = 16'h3d9c;
mem_array[20781] = 16'hebd2;
mem_array[20780] = 16'hbcc4;
mem_array[20783] = 16'h7e31;
mem_array[20782] = 16'hbdd1;
mem_array[20785] = 16'h6a1c;
mem_array[20784] = 16'h3e3d;
mem_array[20787] = 16'hfbdc;
mem_array[20786] = 16'hbf73;
mem_array[20789] = 16'hdc64;
mem_array[20788] = 16'hbd3d;
mem_array[20791] = 16'h5d15;
mem_array[20790] = 16'hbe42;
mem_array[20793] = 16'h36fe;
mem_array[20792] = 16'hbe38;
mem_array[20795] = 16'h55e2;
mem_array[20794] = 16'h3dfb;
mem_array[20797] = 16'h627f;
mem_array[20796] = 16'hbd7b;
mem_array[20799] = 16'h5431;
mem_array[20798] = 16'hbdc9;
mem_array[20801] = 16'h1eda;
mem_array[20800] = 16'h3e79;
mem_array[20803] = 16'hf2a5;
mem_array[20802] = 16'h3e10;
mem_array[20805] = 16'h2aa7;
mem_array[20804] = 16'hbe60;
mem_array[20807] = 16'hac59;
mem_array[20806] = 16'h3c08;
mem_array[20809] = 16'h8e0c;
mem_array[20808] = 16'hbf8f;
mem_array[20811] = 16'h8418;
mem_array[20810] = 16'hbe09;
mem_array[20813] = 16'h0bb4;
mem_array[20812] = 16'h3db0;
mem_array[20815] = 16'h45f0;
mem_array[20814] = 16'h3e32;
mem_array[20817] = 16'h10ab;
mem_array[20816] = 16'hbe92;
mem_array[20819] = 16'hea6d;
mem_array[20818] = 16'h3dec;
mem_array[20821] = 16'hd579;
mem_array[20820] = 16'hbf32;
mem_array[20823] = 16'h4033;
mem_array[20822] = 16'h3e8e;
mem_array[20825] = 16'h930d;
mem_array[20824] = 16'hbf41;
mem_array[20827] = 16'h4815;
mem_array[20826] = 16'h3e95;
mem_array[20829] = 16'he022;
mem_array[20828] = 16'hbe0f;
mem_array[20831] = 16'hc8f5;
mem_array[20830] = 16'h3e2f;
mem_array[20833] = 16'hfb11;
mem_array[20832] = 16'h3e75;
mem_array[20835] = 16'he38a;
mem_array[20834] = 16'h39ee;
mem_array[20837] = 16'h5a3e;
mem_array[20836] = 16'hbed1;
mem_array[20839] = 16'h72b5;
mem_array[20838] = 16'hbeba;
mem_array[20841] = 16'h1811;
mem_array[20840] = 16'hbc43;
mem_array[20843] = 16'h391f;
mem_array[20842] = 16'h3d65;
mem_array[20845] = 16'ha85b;
mem_array[20844] = 16'hba0f;
mem_array[20847] = 16'he522;
mem_array[20846] = 16'hbf8e;
mem_array[20849] = 16'hb1bc;
mem_array[20848] = 16'hbee1;
mem_array[20851] = 16'h70e7;
mem_array[20850] = 16'hbe3c;
mem_array[20853] = 16'haf11;
mem_array[20852] = 16'h3a1b;
mem_array[20855] = 16'h03b2;
mem_array[20854] = 16'h3ec4;
mem_array[20857] = 16'h05b9;
mem_array[20856] = 16'h3e3b;
mem_array[20859] = 16'hee7c;
mem_array[20858] = 16'h3dc0;
mem_array[20861] = 16'h6f76;
mem_array[20860] = 16'h3e89;
mem_array[20863] = 16'hfc99;
mem_array[20862] = 16'hbd66;
mem_array[20865] = 16'hf937;
mem_array[20864] = 16'h3d41;
mem_array[20867] = 16'hc2ed;
mem_array[20866] = 16'h3e27;
mem_array[20869] = 16'hce14;
mem_array[20868] = 16'h3b80;
mem_array[20871] = 16'hf73b;
mem_array[20870] = 16'h3e1f;
mem_array[20873] = 16'hfae8;
mem_array[20872] = 16'h3d99;
mem_array[20875] = 16'h5394;
mem_array[20874] = 16'h3d78;
mem_array[20877] = 16'h4546;
mem_array[20876] = 16'hbd2b;
mem_array[20879] = 16'hbe2a;
mem_array[20878] = 16'h3e56;
mem_array[20881] = 16'h06c7;
mem_array[20880] = 16'hbd49;
mem_array[20883] = 16'haecc;
mem_array[20882] = 16'h3e0f;
mem_array[20885] = 16'h0d34;
mem_array[20884] = 16'hc022;
mem_array[20887] = 16'h8f80;
mem_array[20886] = 16'hbd0a;
mem_array[20889] = 16'h8f0e;
mem_array[20888] = 16'hbe65;
mem_array[20891] = 16'h2208;
mem_array[20890] = 16'h3e82;
mem_array[20893] = 16'h1e7b;
mem_array[20892] = 16'h3e8c;
mem_array[20895] = 16'hd90f;
mem_array[20894] = 16'h3e0e;
mem_array[20897] = 16'hc9b0;
mem_array[20896] = 16'hbdfb;
mem_array[20899] = 16'hebb0;
mem_array[20898] = 16'h3d01;
mem_array[20901] = 16'h1759;
mem_array[20900] = 16'hbc35;
mem_array[20903] = 16'h5470;
mem_array[20902] = 16'h3bac;
mem_array[20905] = 16'hd196;
mem_array[20904] = 16'hbe86;
mem_array[20907] = 16'hc752;
mem_array[20906] = 16'hbf33;
mem_array[20909] = 16'h3447;
mem_array[20908] = 16'hbf43;
mem_array[20911] = 16'h99a1;
mem_array[20910] = 16'h3c62;
mem_array[20913] = 16'h3352;
mem_array[20912] = 16'hbf06;
mem_array[20915] = 16'h4a97;
mem_array[20914] = 16'h3ec9;
mem_array[20917] = 16'h700a;
mem_array[20916] = 16'hbdf0;
mem_array[20919] = 16'hb2eb;
mem_array[20918] = 16'h3d7e;
mem_array[20921] = 16'h622f;
mem_array[20920] = 16'h3ed4;
mem_array[20923] = 16'hd149;
mem_array[20922] = 16'hbd8d;
mem_array[20925] = 16'h7b26;
mem_array[20924] = 16'hbd3d;
mem_array[20927] = 16'h2dd8;
mem_array[20926] = 16'hbc57;
mem_array[20929] = 16'h6b98;
mem_array[20928] = 16'h3e5b;
mem_array[20931] = 16'ha89f;
mem_array[20930] = 16'hbed7;
mem_array[20933] = 16'haabc;
mem_array[20932] = 16'h3d87;
mem_array[20935] = 16'he891;
mem_array[20934] = 16'hbe24;
mem_array[20937] = 16'h7443;
mem_array[20936] = 16'h3e2d;
mem_array[20939] = 16'h3a32;
mem_array[20938] = 16'h3ebe;
mem_array[20941] = 16'hc0fa;
mem_array[20940] = 16'h3d88;
mem_array[20943] = 16'h0d78;
mem_array[20942] = 16'hbf23;
mem_array[20945] = 16'ha641;
mem_array[20944] = 16'hbf9f;
mem_array[20947] = 16'h2d57;
mem_array[20946] = 16'hbe98;
mem_array[20949] = 16'hea8c;
mem_array[20948] = 16'hbe2b;
mem_array[20951] = 16'h99a6;
mem_array[20950] = 16'h3ea3;
mem_array[20953] = 16'hb172;
mem_array[20952] = 16'hbd01;
mem_array[20955] = 16'hfa83;
mem_array[20954] = 16'h3e87;
mem_array[20957] = 16'h226b;
mem_array[20956] = 16'hbea4;
mem_array[20959] = 16'h9534;
mem_array[20958] = 16'h3e58;
mem_array[20961] = 16'hbac9;
mem_array[20960] = 16'hbe06;
mem_array[20963] = 16'hb9a1;
mem_array[20962] = 16'h3ca5;
mem_array[20965] = 16'h90ba;
mem_array[20964] = 16'h3c3d;
mem_array[20967] = 16'hcedb;
mem_array[20966] = 16'hbf10;
mem_array[20969] = 16'h1cad;
mem_array[20968] = 16'hbf6f;
mem_array[20971] = 16'hc5d0;
mem_array[20970] = 16'h3cc3;
mem_array[20973] = 16'hd9f9;
mem_array[20972] = 16'hbee8;
mem_array[20975] = 16'h708c;
mem_array[20974] = 16'hbf0b;
mem_array[20977] = 16'h3323;
mem_array[20976] = 16'hbf2c;
mem_array[20979] = 16'hb50e;
mem_array[20978] = 16'hbdb9;
mem_array[20981] = 16'h1c7b;
mem_array[20980] = 16'h3eac;
mem_array[20983] = 16'h0b8d;
mem_array[20982] = 16'hbde5;
mem_array[20985] = 16'hbe8a;
mem_array[20984] = 16'h3e1b;
mem_array[20987] = 16'h1275;
mem_array[20986] = 16'hbe08;
mem_array[20989] = 16'h6540;
mem_array[20988] = 16'h3e95;
mem_array[20991] = 16'habc0;
mem_array[20990] = 16'hbfc6;
mem_array[20993] = 16'h9df8;
mem_array[20992] = 16'h3e08;
mem_array[20995] = 16'h2004;
mem_array[20994] = 16'hbe17;
mem_array[20997] = 16'h886b;
mem_array[20996] = 16'h3ded;
mem_array[20999] = 16'ha732;
mem_array[20998] = 16'h3e00;
mem_array[21001] = 16'hc3a9;
mem_array[21000] = 16'h3e9f;
mem_array[21003] = 16'h68bb;
mem_array[21002] = 16'hbeba;
mem_array[21005] = 16'h26f7;
mem_array[21004] = 16'hbeb8;
mem_array[21007] = 16'h5a6e;
mem_array[21006] = 16'hbf5d;
mem_array[21009] = 16'hf747;
mem_array[21008] = 16'hbec2;
mem_array[21011] = 16'h1e91;
mem_array[21010] = 16'h3e7b;
mem_array[21013] = 16'h4dd5;
mem_array[21012] = 16'h3e37;
mem_array[21015] = 16'h2b23;
mem_array[21014] = 16'h3e97;
mem_array[21017] = 16'haf4f;
mem_array[21016] = 16'hbd0e;
mem_array[21019] = 16'h523a;
mem_array[21018] = 16'h3d4a;
mem_array[21021] = 16'hcb9d;
mem_array[21020] = 16'hbdd6;
mem_array[21023] = 16'h608d;
mem_array[21022] = 16'h3c96;
mem_array[21025] = 16'h1892;
mem_array[21024] = 16'hbd9f;
mem_array[21027] = 16'hf62c;
mem_array[21026] = 16'hbe84;
mem_array[21029] = 16'h64a9;
mem_array[21028] = 16'hbf42;
mem_array[21031] = 16'hda35;
mem_array[21030] = 16'h3e55;
mem_array[21033] = 16'h6281;
mem_array[21032] = 16'hbe97;
mem_array[21035] = 16'hc456;
mem_array[21034] = 16'hbef7;
mem_array[21037] = 16'h48c1;
mem_array[21036] = 16'hbe33;
mem_array[21039] = 16'h58ab;
mem_array[21038] = 16'hbf35;
mem_array[21041] = 16'he1e7;
mem_array[21040] = 16'h3d82;
mem_array[21043] = 16'h1a68;
mem_array[21042] = 16'h3b84;
mem_array[21045] = 16'h042f;
mem_array[21044] = 16'hbdf0;
mem_array[21047] = 16'h463f;
mem_array[21046] = 16'hbe9b;
mem_array[21049] = 16'h3f7d;
mem_array[21048] = 16'h3ea6;
mem_array[21051] = 16'hc9f5;
mem_array[21050] = 16'hbe57;
mem_array[21053] = 16'h6262;
mem_array[21052] = 16'h3db4;
mem_array[21055] = 16'hd1cd;
mem_array[21054] = 16'hbf20;
mem_array[21057] = 16'h1583;
mem_array[21056] = 16'h3d9a;
mem_array[21059] = 16'hace7;
mem_array[21058] = 16'hbe81;
mem_array[21061] = 16'h3d9c;
mem_array[21060] = 16'h3e57;
mem_array[21063] = 16'h4ba3;
mem_array[21062] = 16'hbf41;
mem_array[21065] = 16'ha18c;
mem_array[21064] = 16'hbe9e;
mem_array[21067] = 16'h5890;
mem_array[21066] = 16'hbf8c;
mem_array[21069] = 16'h38e1;
mem_array[21068] = 16'h3a8a;
mem_array[21071] = 16'hff26;
mem_array[21070] = 16'h3e80;
mem_array[21073] = 16'h1201;
mem_array[21072] = 16'hbd54;
mem_array[21075] = 16'ha24e;
mem_array[21074] = 16'h3e91;
mem_array[21077] = 16'he2d3;
mem_array[21076] = 16'hbe80;
mem_array[21079] = 16'h9b53;
mem_array[21078] = 16'hbb71;
mem_array[21081] = 16'h3c39;
mem_array[21080] = 16'hbd10;
mem_array[21083] = 16'hbf1b;
mem_array[21082] = 16'hbd25;
mem_array[21085] = 16'h9fe2;
mem_array[21084] = 16'hbeea;
mem_array[21087] = 16'h24a2;
mem_array[21086] = 16'hbf4c;
mem_array[21089] = 16'h5ec5;
mem_array[21088] = 16'hbf13;
mem_array[21091] = 16'h8c2b;
mem_array[21090] = 16'h3e89;
mem_array[21093] = 16'h5944;
mem_array[21092] = 16'hbd83;
mem_array[21095] = 16'hed3d;
mem_array[21094] = 16'h3ceb;
mem_array[21097] = 16'h2582;
mem_array[21096] = 16'h3f0e;
mem_array[21099] = 16'hc87b;
mem_array[21098] = 16'hbf42;
mem_array[21101] = 16'h8fe6;
mem_array[21100] = 16'h3e58;
mem_array[21103] = 16'h4061;
mem_array[21102] = 16'h3ec4;
mem_array[21105] = 16'h5f1d;
mem_array[21104] = 16'hbe2f;
mem_array[21107] = 16'hf2fb;
mem_array[21106] = 16'hbe4c;
mem_array[21109] = 16'hd86d;
mem_array[21108] = 16'h3e52;
mem_array[21111] = 16'h2fb1;
mem_array[21110] = 16'h3e43;
mem_array[21113] = 16'hef96;
mem_array[21112] = 16'h3cbb;
mem_array[21115] = 16'ha8e7;
mem_array[21114] = 16'hbf22;
mem_array[21117] = 16'h3a7f;
mem_array[21116] = 16'hbe9a;
mem_array[21119] = 16'h8497;
mem_array[21118] = 16'hbe1a;
mem_array[21121] = 16'hb95b;
mem_array[21120] = 16'h3e8a;
mem_array[21123] = 16'hc14b;
mem_array[21122] = 16'h3e18;
mem_array[21125] = 16'h9229;
mem_array[21124] = 16'hbca4;
mem_array[21127] = 16'h5b6b;
mem_array[21126] = 16'hbf65;
mem_array[21129] = 16'hfd50;
mem_array[21128] = 16'h3e08;
mem_array[21131] = 16'h7893;
mem_array[21130] = 16'h3dc1;
mem_array[21133] = 16'h5d3b;
mem_array[21132] = 16'hbe94;
mem_array[21135] = 16'h075c;
mem_array[21134] = 16'h3e69;
mem_array[21137] = 16'h17a1;
mem_array[21136] = 16'hbdc7;
mem_array[21139] = 16'h6d3d;
mem_array[21138] = 16'h3e18;
mem_array[21141] = 16'h2561;
mem_array[21140] = 16'hbdca;
mem_array[21143] = 16'h0331;
mem_array[21142] = 16'hbc90;
mem_array[21145] = 16'he80e;
mem_array[21144] = 16'hbe7c;
mem_array[21147] = 16'hb872;
mem_array[21146] = 16'hbdfe;
mem_array[21149] = 16'hc392;
mem_array[21148] = 16'hbeba;
mem_array[21151] = 16'h08f3;
mem_array[21150] = 16'h3d15;
mem_array[21153] = 16'h65bc;
mem_array[21152] = 16'h3e89;
mem_array[21155] = 16'h97c3;
mem_array[21154] = 16'h3dae;
mem_array[21157] = 16'he753;
mem_array[21156] = 16'h3e79;
mem_array[21159] = 16'hc041;
mem_array[21158] = 16'hbe9c;
mem_array[21161] = 16'h2dca;
mem_array[21160] = 16'h3e30;
mem_array[21163] = 16'h079a;
mem_array[21162] = 16'hbda6;
mem_array[21165] = 16'hb0d6;
mem_array[21164] = 16'hbea5;
mem_array[21167] = 16'hdb2b;
mem_array[21166] = 16'hbe32;
mem_array[21169] = 16'h6cc6;
mem_array[21168] = 16'h3eae;
mem_array[21171] = 16'h317e;
mem_array[21170] = 16'h3df4;
mem_array[21173] = 16'h2539;
mem_array[21172] = 16'h3d8b;
mem_array[21175] = 16'h5c19;
mem_array[21174] = 16'hbfc6;
mem_array[21177] = 16'hd26b;
mem_array[21176] = 16'h3d91;
mem_array[21179] = 16'hc83d;
mem_array[21178] = 16'hbdca;
mem_array[21181] = 16'h7d07;
mem_array[21180] = 16'h3dee;
mem_array[21183] = 16'h6ce5;
mem_array[21182] = 16'hbcdc;
mem_array[21185] = 16'h99d7;
mem_array[21184] = 16'hbd16;
mem_array[21187] = 16'hb775;
mem_array[21186] = 16'hbf3e;
mem_array[21189] = 16'hbf4b;
mem_array[21188] = 16'h3e58;
mem_array[21191] = 16'h50c8;
mem_array[21190] = 16'hbe2f;
mem_array[21193] = 16'h07ca;
mem_array[21192] = 16'hbe0d;
mem_array[21195] = 16'h726b;
mem_array[21194] = 16'h3ea2;
mem_array[21197] = 16'h69b4;
mem_array[21196] = 16'h3c3f;
mem_array[21199] = 16'hebc7;
mem_array[21198] = 16'hbe3f;
mem_array[21201] = 16'h189e;
mem_array[21200] = 16'hbdb1;
mem_array[21203] = 16'hdd31;
mem_array[21202] = 16'h3d8b;
mem_array[21205] = 16'h5935;
mem_array[21204] = 16'h3e94;
mem_array[21207] = 16'hf373;
mem_array[21206] = 16'hbe7b;
mem_array[21209] = 16'h055e;
mem_array[21208] = 16'hbec6;
mem_array[21211] = 16'h8f0c;
mem_array[21210] = 16'h3e22;
mem_array[21213] = 16'h795d;
mem_array[21212] = 16'h3e07;
mem_array[21215] = 16'hff62;
mem_array[21214] = 16'hbda4;
mem_array[21217] = 16'h3ae7;
mem_array[21216] = 16'h3e73;
mem_array[21219] = 16'h6868;
mem_array[21218] = 16'h3e49;
mem_array[21221] = 16'h3edc;
mem_array[21220] = 16'h3d3d;
mem_array[21223] = 16'h064f;
mem_array[21222] = 16'h3dbb;
mem_array[21225] = 16'h1c22;
mem_array[21224] = 16'h3e93;
mem_array[21227] = 16'h261b;
mem_array[21226] = 16'hbd37;
mem_array[21229] = 16'hc9f1;
mem_array[21228] = 16'hbc6f;
mem_array[21231] = 16'h5f4e;
mem_array[21230] = 16'hbede;
mem_array[21233] = 16'h77db;
mem_array[21232] = 16'h3cb8;
mem_array[21235] = 16'h5935;
mem_array[21234] = 16'hbfd1;
mem_array[21237] = 16'h5241;
mem_array[21236] = 16'hbea0;
mem_array[21239] = 16'h9b40;
mem_array[21238] = 16'h3e07;
mem_array[21241] = 16'h18ae;
mem_array[21240] = 16'hbe69;
mem_array[21243] = 16'h9f9b;
mem_array[21242] = 16'h3e1a;
mem_array[21245] = 16'hc5a3;
mem_array[21244] = 16'hbe52;
mem_array[21247] = 16'h2df9;
mem_array[21246] = 16'h3d70;
mem_array[21249] = 16'hca31;
mem_array[21248] = 16'h3e37;
mem_array[21251] = 16'he6e3;
mem_array[21250] = 16'hbd2a;
mem_array[21253] = 16'hf724;
mem_array[21252] = 16'hbe1a;
mem_array[21255] = 16'h105d;
mem_array[21254] = 16'h3eb0;
mem_array[21257] = 16'hc348;
mem_array[21256] = 16'h3e72;
mem_array[21259] = 16'h2619;
mem_array[21258] = 16'hbed9;
mem_array[21261] = 16'hb2ea;
mem_array[21260] = 16'hbd0e;
mem_array[21263] = 16'he6fc;
mem_array[21262] = 16'h3d84;
mem_array[21265] = 16'hc102;
mem_array[21264] = 16'hbe2c;
mem_array[21267] = 16'h676d;
mem_array[21266] = 16'hbe9c;
mem_array[21269] = 16'h5a1f;
mem_array[21268] = 16'hbeab;
mem_array[21271] = 16'hcbd3;
mem_array[21270] = 16'h3db0;
mem_array[21273] = 16'hce8c;
mem_array[21272] = 16'h3e2f;
mem_array[21275] = 16'hefb4;
mem_array[21274] = 16'h3e0d;
mem_array[21277] = 16'h9619;
mem_array[21276] = 16'h3e6d;
mem_array[21279] = 16'h2db8;
mem_array[21278] = 16'h3e24;
mem_array[21281] = 16'h4a13;
mem_array[21280] = 16'hbdc9;
mem_array[21283] = 16'h4bfd;
mem_array[21282] = 16'h3e4a;
mem_array[21285] = 16'hdbdd;
mem_array[21284] = 16'h3dee;
mem_array[21287] = 16'hef47;
mem_array[21286] = 16'hbe9a;
mem_array[21289] = 16'h5421;
mem_array[21288] = 16'h3e14;
mem_array[21291] = 16'h771a;
mem_array[21290] = 16'hbe36;
mem_array[21293] = 16'h11a8;
mem_array[21292] = 16'hbd59;
mem_array[21295] = 16'h043f;
mem_array[21294] = 16'hc003;
mem_array[21297] = 16'he248;
mem_array[21296] = 16'hbdcd;
mem_array[21299] = 16'hd899;
mem_array[21298] = 16'h3d0b;
mem_array[21301] = 16'h66df;
mem_array[21300] = 16'hbe98;
mem_array[21303] = 16'he811;
mem_array[21302] = 16'hbe5c;
mem_array[21305] = 16'h1eb5;
mem_array[21304] = 16'h3976;
mem_array[21307] = 16'hb52c;
mem_array[21306] = 16'h3e40;
mem_array[21309] = 16'h0957;
mem_array[21308] = 16'h3de7;
mem_array[21311] = 16'hd45b;
mem_array[21310] = 16'hbf38;
mem_array[21313] = 16'hef09;
mem_array[21312] = 16'hbf14;
mem_array[21315] = 16'h1035;
mem_array[21314] = 16'hbd97;
mem_array[21317] = 16'h778d;
mem_array[21316] = 16'hbe3d;
mem_array[21319] = 16'h8c5e;
mem_array[21318] = 16'hbf84;
mem_array[21321] = 16'hbaa9;
mem_array[21320] = 16'hbe2f;
mem_array[21323] = 16'hdc17;
mem_array[21322] = 16'hbd6f;
mem_array[21325] = 16'h0c7e;
mem_array[21324] = 16'h3df9;
mem_array[21327] = 16'h4999;
mem_array[21326] = 16'hbd18;
mem_array[21329] = 16'h0836;
mem_array[21328] = 16'hbefb;
mem_array[21331] = 16'h89b5;
mem_array[21330] = 16'h3e4c;
mem_array[21333] = 16'he2e9;
mem_array[21332] = 16'h3dac;
mem_array[21335] = 16'hb47b;
mem_array[21334] = 16'hbd0b;
mem_array[21337] = 16'hb12a;
mem_array[21336] = 16'h3c51;
mem_array[21339] = 16'h3002;
mem_array[21338] = 16'h3d88;
mem_array[21341] = 16'he536;
mem_array[21340] = 16'hbdc6;
mem_array[21343] = 16'h618a;
mem_array[21342] = 16'hbdc1;
mem_array[21345] = 16'hf18a;
mem_array[21344] = 16'hbf09;
mem_array[21347] = 16'hb3b0;
mem_array[21346] = 16'hbe16;
mem_array[21349] = 16'h9f79;
mem_array[21348] = 16'hbe58;
mem_array[21351] = 16'h686e;
mem_array[21350] = 16'hbde3;
mem_array[21353] = 16'h7c5d;
mem_array[21352] = 16'hbdee;
mem_array[21355] = 16'ha583;
mem_array[21354] = 16'hc015;
mem_array[21357] = 16'hbe14;
mem_array[21356] = 16'hbea3;
mem_array[21359] = 16'h8f12;
mem_array[21358] = 16'hbef0;
mem_array[21361] = 16'hf496;
mem_array[21360] = 16'hbf10;
mem_array[21363] = 16'h6d0b;
mem_array[21362] = 16'h3dea;
mem_array[21365] = 16'h9d17;
mem_array[21364] = 16'hbe08;
mem_array[21367] = 16'h727d;
mem_array[21366] = 16'hbe0d;
mem_array[21369] = 16'h351b;
mem_array[21368] = 16'hbdf2;
mem_array[21371] = 16'hc6ba;
mem_array[21370] = 16'hbf44;
mem_array[21373] = 16'h2ee5;
mem_array[21372] = 16'hbdc0;
mem_array[21375] = 16'h57fb;
mem_array[21374] = 16'h3e46;
mem_array[21377] = 16'h9dbf;
mem_array[21376] = 16'h3dff;
mem_array[21379] = 16'hec99;
mem_array[21378] = 16'h3e14;
mem_array[21381] = 16'he065;
mem_array[21380] = 16'hbe01;
mem_array[21383] = 16'h924b;
mem_array[21382] = 16'hbc15;
mem_array[21385] = 16'h793c;
mem_array[21384] = 16'hbc80;
mem_array[21387] = 16'h36f2;
mem_array[21386] = 16'h3dc8;
mem_array[21389] = 16'h5c81;
mem_array[21388] = 16'h3ce4;
mem_array[21391] = 16'h9763;
mem_array[21390] = 16'h3e04;
mem_array[21393] = 16'h13e0;
mem_array[21392] = 16'hbee5;
mem_array[21395] = 16'he397;
mem_array[21394] = 16'hbea2;
mem_array[21397] = 16'h94ce;
mem_array[21396] = 16'hbd9a;
mem_array[21399] = 16'h8e3e;
mem_array[21398] = 16'h3c39;
mem_array[21401] = 16'hc3dc;
mem_array[21400] = 16'h3cbc;
mem_array[21403] = 16'h8712;
mem_array[21402] = 16'hbc31;
mem_array[21405] = 16'heaef;
mem_array[21404] = 16'hbe96;
mem_array[21407] = 16'he02d;
mem_array[21406] = 16'h3d81;
mem_array[21409] = 16'he2da;
mem_array[21408] = 16'hbdcb;
mem_array[21411] = 16'hdde8;
mem_array[21410] = 16'hbe44;
mem_array[21413] = 16'h3f95;
mem_array[21412] = 16'hbca7;
mem_array[21415] = 16'h785a;
mem_array[21414] = 16'hbfbc;
mem_array[21417] = 16'h83c4;
mem_array[21416] = 16'hbe97;
mem_array[21419] = 16'heb37;
mem_array[21418] = 16'hbeb9;
mem_array[21421] = 16'h45cf;
mem_array[21420] = 16'h3ec6;
mem_array[21423] = 16'h8d0c;
mem_array[21422] = 16'h3e1e;
mem_array[21425] = 16'hb0ad;
mem_array[21424] = 16'h3bc4;
mem_array[21427] = 16'hfbed;
mem_array[21426] = 16'h3e75;
mem_array[21429] = 16'h6e53;
mem_array[21428] = 16'h3cbb;
mem_array[21431] = 16'hdafc;
mem_array[21430] = 16'hbfa2;
mem_array[21433] = 16'h066c;
mem_array[21432] = 16'hbe54;
mem_array[21435] = 16'h8695;
mem_array[21434] = 16'h3e98;
mem_array[21437] = 16'h895f;
mem_array[21436] = 16'h3e2a;
mem_array[21439] = 16'hab1e;
mem_array[21438] = 16'hbd9e;
mem_array[21441] = 16'h8a14;
mem_array[21440] = 16'hbe0e;
mem_array[21443] = 16'h0276;
mem_array[21442] = 16'h3d5c;
mem_array[21445] = 16'h7e9f;
mem_array[21444] = 16'h3e08;
mem_array[21447] = 16'h2fa2;
mem_array[21446] = 16'h3e06;
mem_array[21449] = 16'h4511;
mem_array[21448] = 16'hbda2;
mem_array[21451] = 16'h2ced;
mem_array[21450] = 16'h3d54;
mem_array[21453] = 16'h31e3;
mem_array[21452] = 16'hbf20;
mem_array[21455] = 16'h5089;
mem_array[21454] = 16'h3dbf;
mem_array[21457] = 16'he2e6;
mem_array[21456] = 16'h3db7;
mem_array[21459] = 16'h972f;
mem_array[21458] = 16'hbd05;
mem_array[21461] = 16'h4bd8;
mem_array[21460] = 16'h3c0e;
mem_array[21463] = 16'h1535;
mem_array[21462] = 16'hbe45;
mem_array[21465] = 16'hf785;
mem_array[21464] = 16'hbeab;
mem_array[21467] = 16'hbeae;
mem_array[21466] = 16'h3c42;
mem_array[21469] = 16'h56fa;
mem_array[21468] = 16'hbe9f;
mem_array[21471] = 16'h6ca4;
mem_array[21470] = 16'hbec0;
mem_array[21473] = 16'h54e4;
mem_array[21472] = 16'hbdb8;
mem_array[21475] = 16'hbf55;
mem_array[21474] = 16'hbf69;
mem_array[21477] = 16'hacef;
mem_array[21476] = 16'hbe1d;
mem_array[21479] = 16'hb984;
mem_array[21478] = 16'hbefb;
mem_array[21481] = 16'h112f;
mem_array[21480] = 16'h3dc6;
mem_array[21483] = 16'h4ae3;
mem_array[21482] = 16'hbe0f;
mem_array[21485] = 16'h25a6;
mem_array[21484] = 16'hbb63;
mem_array[21487] = 16'hfdfc;
mem_array[21486] = 16'h3e54;
mem_array[21489] = 16'ha10e;
mem_array[21488] = 16'h3e94;
mem_array[21491] = 16'h7582;
mem_array[21490] = 16'hbf7a;
mem_array[21493] = 16'h8da4;
mem_array[21492] = 16'hbf62;
mem_array[21495] = 16'hf273;
mem_array[21494] = 16'hbde3;
mem_array[21497] = 16'h7f0f;
mem_array[21496] = 16'h3d78;
mem_array[21499] = 16'h480b;
mem_array[21498] = 16'h3ea2;
mem_array[21501] = 16'h9a98;
mem_array[21500] = 16'hbd26;
mem_array[21503] = 16'ha08b;
mem_array[21502] = 16'hbd60;
mem_array[21505] = 16'hab2d;
mem_array[21504] = 16'h3c68;
mem_array[21507] = 16'ha737;
mem_array[21506] = 16'h3db6;
mem_array[21509] = 16'h5278;
mem_array[21508] = 16'h3db3;
mem_array[21511] = 16'h276a;
mem_array[21510] = 16'h3edb;
mem_array[21513] = 16'he6fb;
mem_array[21512] = 16'hbfb2;
mem_array[21515] = 16'h5be1;
mem_array[21514] = 16'h3ea8;
mem_array[21517] = 16'h02ae;
mem_array[21516] = 16'h3e9b;
mem_array[21519] = 16'hf45c;
mem_array[21518] = 16'hbd3f;
mem_array[21521] = 16'hfbc7;
mem_array[21520] = 16'hbd80;
mem_array[21523] = 16'hab44;
mem_array[21522] = 16'hbd88;
mem_array[21525] = 16'hb0b4;
mem_array[21524] = 16'hbf13;
mem_array[21527] = 16'hdcbb;
mem_array[21526] = 16'h3e92;
mem_array[21529] = 16'h1f5d;
mem_array[21528] = 16'hbf16;
mem_array[21531] = 16'hef57;
mem_array[21530] = 16'hbe62;
mem_array[21533] = 16'h4bcf;
mem_array[21532] = 16'hbf02;
mem_array[21535] = 16'ha31c;
mem_array[21534] = 16'hbf20;
mem_array[21537] = 16'h82e1;
mem_array[21536] = 16'hbe86;
mem_array[21539] = 16'h31bc;
mem_array[21538] = 16'hbf23;
mem_array[21541] = 16'h1ced;
mem_array[21540] = 16'hbf20;
mem_array[21543] = 16'hd605;
mem_array[21542] = 16'hbdcb;
mem_array[21545] = 16'hcde9;
mem_array[21544] = 16'hbef8;
mem_array[21547] = 16'h5874;
mem_array[21546] = 16'h3f01;
mem_array[21549] = 16'hb3d8;
mem_array[21548] = 16'hbd02;
mem_array[21551] = 16'hd452;
mem_array[21550] = 16'hbf2c;
mem_array[21553] = 16'h71fb;
mem_array[21552] = 16'hbe80;
mem_array[21555] = 16'h16ad;
mem_array[21554] = 16'hbeb5;
mem_array[21557] = 16'h0f6a;
mem_array[21556] = 16'hbea7;
mem_array[21559] = 16'hc839;
mem_array[21558] = 16'h3ee0;
mem_array[21561] = 16'h264f;
mem_array[21560] = 16'hbc93;
mem_array[21563] = 16'hacef;
mem_array[21562] = 16'h3ca3;
mem_array[21565] = 16'h43db;
mem_array[21564] = 16'hbd43;
mem_array[21567] = 16'h3ad8;
mem_array[21566] = 16'hbe56;
mem_array[21569] = 16'hec73;
mem_array[21568] = 16'hbea5;
mem_array[21571] = 16'hdcca;
mem_array[21570] = 16'h3f3b;
mem_array[21573] = 16'hafb5;
mem_array[21572] = 16'hbf40;
mem_array[21575] = 16'h8151;
mem_array[21574] = 16'hbe4c;
mem_array[21577] = 16'h5b14;
mem_array[21576] = 16'h3edc;
mem_array[21579] = 16'h5d80;
mem_array[21578] = 16'hbf06;
mem_array[21581] = 16'h7c48;
mem_array[21580] = 16'h3e01;
mem_array[21583] = 16'h9019;
mem_array[21582] = 16'hbe19;
mem_array[21585] = 16'h3942;
mem_array[21584] = 16'hbe52;
mem_array[21587] = 16'hc8b3;
mem_array[21586] = 16'h3ee3;
mem_array[21589] = 16'h5efe;
mem_array[21588] = 16'hbdd4;
mem_array[21591] = 16'h1d85;
mem_array[21590] = 16'hbf7e;
mem_array[21593] = 16'hc992;
mem_array[21592] = 16'hbe8d;
mem_array[21595] = 16'h68b5;
mem_array[21594] = 16'hbf21;
mem_array[21597] = 16'hab6f;
mem_array[21596] = 16'hbe9a;
mem_array[21599] = 16'h911e;
mem_array[21598] = 16'hbecf;
mem_array[21601] = 16'h0987;
mem_array[21600] = 16'hbedc;
mem_array[21603] = 16'h8610;
mem_array[21602] = 16'hbe9e;
mem_array[21605] = 16'h85db;
mem_array[21604] = 16'hbce6;
mem_array[21607] = 16'h15be;
mem_array[21606] = 16'h3eb8;
mem_array[21609] = 16'h7892;
mem_array[21608] = 16'hbfaa;
mem_array[21611] = 16'h8daf;
mem_array[21610] = 16'h3ae9;
mem_array[21613] = 16'h5cb3;
mem_array[21612] = 16'h3f5c;
mem_array[21615] = 16'h8313;
mem_array[21614] = 16'hbea8;
mem_array[21617] = 16'h90d5;
mem_array[21616] = 16'h3ef3;
mem_array[21619] = 16'he708;
mem_array[21618] = 16'hbe70;
mem_array[21621] = 16'hd889;
mem_array[21620] = 16'h3c40;
mem_array[21623] = 16'haab6;
mem_array[21622] = 16'hbbcf;
mem_array[21625] = 16'he0b5;
mem_array[21624] = 16'h3e11;
mem_array[21627] = 16'hbf39;
mem_array[21626] = 16'h3e64;
mem_array[21629] = 16'hf7e2;
mem_array[21628] = 16'hbe58;
mem_array[21631] = 16'h2dfd;
mem_array[21630] = 16'h3f10;
mem_array[21633] = 16'hc50d;
mem_array[21632] = 16'hbf37;
mem_array[21635] = 16'h34c0;
mem_array[21634] = 16'hbda4;
mem_array[21637] = 16'hb5d0;
mem_array[21636] = 16'hbf6c;
mem_array[21639] = 16'h50e6;
mem_array[21638] = 16'hbf14;
mem_array[21641] = 16'hfaec;
mem_array[21640] = 16'h3da7;
mem_array[21643] = 16'h7382;
mem_array[21642] = 16'h3e57;
mem_array[21645] = 16'he895;
mem_array[21644] = 16'hbf1d;
mem_array[21647] = 16'h2e4e;
mem_array[21646] = 16'h3eb1;
mem_array[21649] = 16'ha696;
mem_array[21648] = 16'hbb3b;
mem_array[21651] = 16'h91dd;
mem_array[21650] = 16'hbf8d;
mem_array[21653] = 16'h0af7;
mem_array[21652] = 16'hbee1;
mem_array[21655] = 16'he3b3;
mem_array[21654] = 16'h3f3d;
mem_array[21657] = 16'he57d;
mem_array[21656] = 16'h3c73;
mem_array[21659] = 16'he247;
mem_array[21658] = 16'hbe5a;
mem_array[21661] = 16'hc10d;
mem_array[21660] = 16'hbe6e;
mem_array[21663] = 16'h270a;
mem_array[21662] = 16'hbf1c;
mem_array[21665] = 16'h1f9e;
mem_array[21664] = 16'h3d88;
mem_array[21667] = 16'h0a7e;
mem_array[21666] = 16'hbeb9;
mem_array[21669] = 16'h47d8;
mem_array[21668] = 16'hbe2f;
mem_array[21671] = 16'h806c;
mem_array[21670] = 16'hbee6;
mem_array[21673] = 16'hc16a;
mem_array[21672] = 16'h3f9f;
mem_array[21675] = 16'hc76a;
mem_array[21674] = 16'h3e93;
mem_array[21677] = 16'h29a7;
mem_array[21676] = 16'h3f79;
mem_array[21679] = 16'h5953;
mem_array[21678] = 16'h3e41;
mem_array[21681] = 16'h360b;
mem_array[21680] = 16'hbd2f;
mem_array[21683] = 16'hf870;
mem_array[21682] = 16'hbcaa;
mem_array[21685] = 16'h8e98;
mem_array[21684] = 16'hbed7;
mem_array[21687] = 16'h1f4f;
mem_array[21686] = 16'h3e50;
mem_array[21689] = 16'h2c60;
mem_array[21688] = 16'h3f06;
mem_array[21691] = 16'h47e8;
mem_array[21690] = 16'h3e02;
mem_array[21693] = 16'h8b54;
mem_array[21692] = 16'hbedd;
mem_array[21695] = 16'hd6db;
mem_array[21694] = 16'h3f5b;
mem_array[21697] = 16'hee6d;
mem_array[21696] = 16'hbe88;
mem_array[21699] = 16'h735e;
mem_array[21698] = 16'h3f47;
mem_array[21701] = 16'hcab9;
mem_array[21700] = 16'h3f18;
mem_array[21703] = 16'h39e1;
mem_array[21702] = 16'h3f08;
mem_array[21705] = 16'h66f1;
mem_array[21704] = 16'hbf51;
mem_array[21707] = 16'h1ea4;
mem_array[21706] = 16'h3d9b;
mem_array[21709] = 16'hb2e3;
mem_array[21708] = 16'h3f89;
mem_array[21711] = 16'hb9cb;
mem_array[21710] = 16'hbd26;
mem_array[21713] = 16'hafcf;
mem_array[21712] = 16'h3ed9;
mem_array[21715] = 16'h0201;
mem_array[21714] = 16'h3f77;
mem_array[21717] = 16'h7f7d;
mem_array[21716] = 16'h3fc1;
mem_array[21719] = 16'h11de;
mem_array[21718] = 16'h3dc2;
mem_array[21721] = 16'h1c8c;
mem_array[21720] = 16'hbf97;
mem_array[21723] = 16'h65bf;
mem_array[21722] = 16'hbea9;
mem_array[21725] = 16'hddd6;
mem_array[21724] = 16'h3ef8;
mem_array[21727] = 16'h6388;
mem_array[21726] = 16'hbf32;
mem_array[21729] = 16'h78d8;
mem_array[21728] = 16'h3eb6;
mem_array[21731] = 16'hbc01;
mem_array[21730] = 16'hbe03;
mem_array[21733] = 16'h680b;
mem_array[21732] = 16'hbf15;
mem_array[21735] = 16'hd514;
mem_array[21734] = 16'h3e98;
mem_array[21737] = 16'hae5a;
mem_array[21736] = 16'hbceb;
mem_array[21739] = 16'hc956;
mem_array[21738] = 16'hbdee;
mem_array[21741] = 16'h0f6c;
mem_array[21740] = 16'h3cd9;
mem_array[21743] = 16'h4e45;
mem_array[21742] = 16'hbcd8;
mem_array[21745] = 16'hebbc;
mem_array[21744] = 16'hbfc7;
mem_array[21747] = 16'hae6a;
mem_array[21746] = 16'h3eda;
mem_array[21749] = 16'h890a;
mem_array[21748] = 16'h3fa8;
mem_array[21751] = 16'hbef1;
mem_array[21750] = 16'h3f37;
mem_array[21753] = 16'he530;
mem_array[21752] = 16'hbed2;
mem_array[21755] = 16'h4190;
mem_array[21754] = 16'hbe29;
mem_array[21757] = 16'h0134;
mem_array[21756] = 16'hbf48;
mem_array[21759] = 16'h43b6;
mem_array[21758] = 16'h3f05;
mem_array[21761] = 16'hd0b1;
mem_array[21760] = 16'h3bbf;
mem_array[21763] = 16'hee35;
mem_array[21762] = 16'h3f28;
mem_array[21765] = 16'had19;
mem_array[21764] = 16'hbf9e;
mem_array[21767] = 16'hd217;
mem_array[21766] = 16'hbf49;
mem_array[21769] = 16'ha948;
mem_array[21768] = 16'h3e72;
mem_array[21771] = 16'hbd23;
mem_array[21770] = 16'hbc7a;
mem_array[21773] = 16'haa46;
mem_array[21772] = 16'h3ed0;
mem_array[21775] = 16'h15b6;
mem_array[21774] = 16'h3f0a;
mem_array[21777] = 16'h3118;
mem_array[21776] = 16'h3fc7;
mem_array[21779] = 16'hdcf5;
mem_array[21778] = 16'hbde1;
mem_array[21781] = 16'h5a16;
mem_array[21780] = 16'h3c8b;
mem_array[21783] = 16'h1b9e;
mem_array[21782] = 16'hbda4;
mem_array[21785] = 16'h85c7;
mem_array[21784] = 16'h3d88;
mem_array[21787] = 16'he1bb;
mem_array[21786] = 16'h3daa;
mem_array[21789] = 16'h0d55;
mem_array[21788] = 16'h3d47;
mem_array[21791] = 16'h77f5;
mem_array[21790] = 16'h3f17;
mem_array[21793] = 16'h6c13;
mem_array[21792] = 16'hbe8c;
mem_array[21795] = 16'h64cd;
mem_array[21794] = 16'h3e7c;
mem_array[21797] = 16'haab5;
mem_array[21796] = 16'h3f6c;
mem_array[21799] = 16'hfc56;
mem_array[21798] = 16'h3f8a;
mem_array[21801] = 16'h9637;
mem_array[21800] = 16'h3d20;
mem_array[21803] = 16'h1f16;
mem_array[21802] = 16'hbc77;
mem_array[21805] = 16'h3496;
mem_array[21804] = 16'h3dc4;
mem_array[21807] = 16'h01e5;
mem_array[21806] = 16'hbe13;
mem_array[21809] = 16'h8331;
mem_array[21808] = 16'h3d00;
mem_array[21811] = 16'hbc23;
mem_array[21810] = 16'h3db0;
mem_array[21813] = 16'h8c0a;
mem_array[21812] = 16'hbdcc;
mem_array[21815] = 16'hcc9e;
mem_array[21814] = 16'hbeb2;
mem_array[21817] = 16'hd9d9;
mem_array[21816] = 16'hbcc3;
mem_array[21819] = 16'h1dd8;
mem_array[21818] = 16'h3d0c;
mem_array[21821] = 16'h563a;
mem_array[21820] = 16'hbe45;
mem_array[21823] = 16'h6c70;
mem_array[21822] = 16'hbef3;
mem_array[21825] = 16'hd3d0;
mem_array[21824] = 16'hbde2;
mem_array[21827] = 16'h668f;
mem_array[21826] = 16'hbf5c;
mem_array[21829] = 16'hba11;
mem_array[21828] = 16'hbf07;
mem_array[21831] = 16'hdd8c;
mem_array[21830] = 16'h3d36;
mem_array[21833] = 16'h0550;
mem_array[21832] = 16'hbe78;
mem_array[21835] = 16'hd175;
mem_array[21834] = 16'h3d3d;
mem_array[21837] = 16'hb221;
mem_array[21836] = 16'h3f05;
mem_array[21839] = 16'h9e95;
mem_array[21838] = 16'hbe87;
mem_array[21841] = 16'hb1f5;
mem_array[21840] = 16'hbdd0;
mem_array[21843] = 16'h0122;
mem_array[21842] = 16'hbc92;
mem_array[21845] = 16'h93a5;
mem_array[21844] = 16'hbd28;
mem_array[21847] = 16'h5655;
mem_array[21846] = 16'h3c5c;
mem_array[21849] = 16'h2530;
mem_array[21848] = 16'hbcb2;
mem_array[21851] = 16'h3cbf;
mem_array[21850] = 16'h3d10;
mem_array[21853] = 16'h79bd;
mem_array[21852] = 16'h3d13;
mem_array[21855] = 16'hce25;
mem_array[21854] = 16'hbcff;
mem_array[21857] = 16'he900;
mem_array[21856] = 16'h3d2e;
mem_array[21859] = 16'h36bf;
mem_array[21858] = 16'hbe02;
mem_array[21861] = 16'h85e1;
mem_array[21860] = 16'h3d57;
mem_array[21863] = 16'h0c9a;
mem_array[21862] = 16'h3d9c;
mem_array[21865] = 16'h1639;
mem_array[21864] = 16'h3ba1;
mem_array[21867] = 16'h0ebb;
mem_array[21866] = 16'h3da3;
mem_array[21869] = 16'h27e2;
mem_array[21868] = 16'hbde7;
mem_array[21871] = 16'hf9fa;
mem_array[21870] = 16'h3da5;
mem_array[21873] = 16'h1106;
mem_array[21872] = 16'h3c0a;
mem_array[21875] = 16'h1a0e;
mem_array[21874] = 16'hbddf;
mem_array[21877] = 16'h4bc9;
mem_array[21876] = 16'h3ca4;
mem_array[21879] = 16'h0055;
mem_array[21878] = 16'hbdd5;
mem_array[21881] = 16'h44aa;
mem_array[21880] = 16'hbc0a;
mem_array[21883] = 16'hf3c9;
mem_array[21882] = 16'hbd65;
mem_array[21885] = 16'h88f8;
mem_array[21884] = 16'hbc2b;
mem_array[21887] = 16'hbd93;
mem_array[21886] = 16'hbd32;
mem_array[21889] = 16'h084e;
mem_array[21888] = 16'h3cb0;
mem_array[21891] = 16'hbbe3;
mem_array[21890] = 16'h3b28;
mem_array[21893] = 16'h1598;
mem_array[21892] = 16'h3cc2;
mem_array[21895] = 16'h6262;
mem_array[21894] = 16'hbdbf;
mem_array[21897] = 16'h8d70;
mem_array[21896] = 16'h3c3e;
mem_array[21899] = 16'h3372;
mem_array[21898] = 16'h3d12;
mem_array[21901] = 16'h863e;
mem_array[21900] = 16'hbbda;
mem_array[21903] = 16'h9089;
mem_array[21902] = 16'hbd6d;
mem_array[21905] = 16'h5c77;
mem_array[21904] = 16'hbddd;
mem_array[21907] = 16'h44cb;
mem_array[21906] = 16'h3e3e;
mem_array[21909] = 16'he74c;
mem_array[21908] = 16'hbd6f;
mem_array[21911] = 16'h1fdb;
mem_array[21910] = 16'hbd15;
mem_array[21913] = 16'he3cc;
mem_array[21912] = 16'hbde4;
mem_array[21915] = 16'h49e5;
mem_array[21914] = 16'h3e79;
mem_array[21917] = 16'hf9ed;
mem_array[21916] = 16'hbd6f;
mem_array[21919] = 16'hadc3;
mem_array[21918] = 16'h3d08;
mem_array[21921] = 16'h8456;
mem_array[21920] = 16'hbccb;
mem_array[21923] = 16'h94aa;
mem_array[21922] = 16'hbdb6;
mem_array[21925] = 16'h2bad;
mem_array[21924] = 16'h3f11;
mem_array[21927] = 16'h4fae;
mem_array[21926] = 16'hbf08;
mem_array[21929] = 16'h9031;
mem_array[21928] = 16'hbd87;
mem_array[21931] = 16'h7e4e;
mem_array[21930] = 16'hbe6b;
mem_array[21933] = 16'h4061;
mem_array[21932] = 16'hbdeb;
mem_array[21935] = 16'h4950;
mem_array[21934] = 16'h3f01;
mem_array[21937] = 16'hbd67;
mem_array[21936] = 16'h3f17;
mem_array[21939] = 16'h4c19;
mem_array[21938] = 16'h3e94;
mem_array[21941] = 16'h947e;
mem_array[21940] = 16'h3d34;
mem_array[21943] = 16'h1d87;
mem_array[21942] = 16'hbe32;
mem_array[21945] = 16'h8e78;
mem_array[21944] = 16'hbd94;
mem_array[21947] = 16'h8c09;
mem_array[21946] = 16'hbdff;
mem_array[21949] = 16'hfbf1;
mem_array[21948] = 16'hbf0c;
mem_array[21951] = 16'h9a67;
mem_array[21950] = 16'h3e00;
mem_array[21953] = 16'hd155;
mem_array[21952] = 16'hbe58;
mem_array[21955] = 16'h5ad5;
mem_array[21954] = 16'h3da0;
mem_array[21957] = 16'hb74a;
mem_array[21956] = 16'hbf0e;
mem_array[21959] = 16'h451e;
mem_array[21958] = 16'hbe51;
mem_array[21961] = 16'he60b;
mem_array[21960] = 16'hbea7;
mem_array[21963] = 16'hd213;
mem_array[21962] = 16'h3f2e;
mem_array[21965] = 16'h75d8;
mem_array[21964] = 16'h3e50;
mem_array[21967] = 16'h4833;
mem_array[21966] = 16'h3e43;
mem_array[21969] = 16'h67e0;
mem_array[21968] = 16'h3cda;
mem_array[21971] = 16'h1787;
mem_array[21970] = 16'hbe6d;
mem_array[21973] = 16'h60cd;
mem_array[21972] = 16'hbf17;
mem_array[21975] = 16'h54fa;
mem_array[21974] = 16'h3d42;
mem_array[21977] = 16'h6626;
mem_array[21976] = 16'h3ee8;
mem_array[21979] = 16'hdca5;
mem_array[21978] = 16'h3d65;
mem_array[21981] = 16'h51ff;
mem_array[21980] = 16'hbda0;
mem_array[21983] = 16'h986e;
mem_array[21982] = 16'hbd12;
mem_array[21985] = 16'hd4a7;
mem_array[21984] = 16'hbf5b;
mem_array[21987] = 16'h4753;
mem_array[21986] = 16'hbeb5;
mem_array[21989] = 16'h4fa2;
mem_array[21988] = 16'h3e86;
mem_array[21991] = 16'hec03;
mem_array[21990] = 16'hbc59;
mem_array[21993] = 16'h494b;
mem_array[21992] = 16'h3eb2;
mem_array[21995] = 16'hda5c;
mem_array[21994] = 16'hbe79;
mem_array[21997] = 16'h6c1f;
mem_array[21996] = 16'h3eda;
mem_array[21999] = 16'h8c78;
mem_array[21998] = 16'hbe2b;
mem_array[22001] = 16'h7884;
mem_array[22000] = 16'hbf64;
mem_array[22003] = 16'hb61e;
mem_array[22002] = 16'h3ebf;
mem_array[22005] = 16'hf15f;
mem_array[22004] = 16'hbdef;
mem_array[22007] = 16'hfacb;
mem_array[22006] = 16'hbf15;
mem_array[22009] = 16'h945c;
mem_array[22008] = 16'hbee5;
mem_array[22011] = 16'he8d4;
mem_array[22010] = 16'h3f72;
mem_array[22013] = 16'h850a;
mem_array[22012] = 16'h3e2e;
mem_array[22015] = 16'hfe70;
mem_array[22014] = 16'h3e8d;
mem_array[22017] = 16'h4cee;
mem_array[22016] = 16'hbf0c;
mem_array[22019] = 16'h79f4;
mem_array[22018] = 16'hbf86;
mem_array[22021] = 16'hc15d;
mem_array[22020] = 16'h3e32;
mem_array[22023] = 16'h37f7;
mem_array[22022] = 16'hbdd2;
mem_array[22025] = 16'hffef;
mem_array[22024] = 16'h3f62;
mem_array[22027] = 16'h230a;
mem_array[22026] = 16'hbf01;
mem_array[22029] = 16'h9c6c;
mem_array[22028] = 16'hbd6f;
mem_array[22031] = 16'h99aa;
mem_array[22030] = 16'hbe28;
mem_array[22033] = 16'hd1dc;
mem_array[22032] = 16'hbcf1;
mem_array[22035] = 16'hd265;
mem_array[22034] = 16'h3fad;
mem_array[22037] = 16'h11f6;
mem_array[22036] = 16'hbf0b;
mem_array[22039] = 16'h8f30;
mem_array[22038] = 16'hbe39;
mem_array[22041] = 16'h8421;
mem_array[22040] = 16'hbd00;
mem_array[22043] = 16'h3906;
mem_array[22042] = 16'h3d5a;
mem_array[22045] = 16'h08aa;
mem_array[22044] = 16'hbfad;
mem_array[22047] = 16'h4d24;
mem_array[22046] = 16'hbf48;
mem_array[22049] = 16'h1c31;
mem_array[22048] = 16'hbf51;
mem_array[22051] = 16'hdd64;
mem_array[22050] = 16'hbdc2;
mem_array[22053] = 16'h7a92;
mem_array[22052] = 16'h3f29;
mem_array[22055] = 16'h33b4;
mem_array[22054] = 16'h3cfb;
mem_array[22057] = 16'hc2fe;
mem_array[22056] = 16'hbd91;
mem_array[22059] = 16'h146d;
mem_array[22058] = 16'hbf0d;
mem_array[22061] = 16'h126f;
mem_array[22060] = 16'hbf43;
mem_array[22063] = 16'h21ea;
mem_array[22062] = 16'hbe19;
mem_array[22065] = 16'had29;
mem_array[22064] = 16'hbf04;
mem_array[22067] = 16'h9505;
mem_array[22066] = 16'h3dd4;
mem_array[22069] = 16'h142d;
mem_array[22068] = 16'hbf80;
mem_array[22071] = 16'h7cff;
mem_array[22070] = 16'h3c73;
mem_array[22073] = 16'h0bc7;
mem_array[22072] = 16'hbedf;
mem_array[22075] = 16'hf07e;
mem_array[22074] = 16'h3d8f;
mem_array[22077] = 16'h240c;
mem_array[22076] = 16'hbe11;
mem_array[22079] = 16'h4ff7;
mem_array[22078] = 16'h3f13;
mem_array[22081] = 16'h8449;
mem_array[22080] = 16'h3e15;
mem_array[22083] = 16'h17b9;
mem_array[22082] = 16'hbee8;
mem_array[22085] = 16'h4458;
mem_array[22084] = 16'hbe4a;
mem_array[22087] = 16'hff0e;
mem_array[22086] = 16'hbccc;
mem_array[22089] = 16'h47c6;
mem_array[22088] = 16'hbe63;
mem_array[22091] = 16'h1786;
mem_array[22090] = 16'h3e35;
mem_array[22093] = 16'h29ba;
mem_array[22092] = 16'h3e95;
mem_array[22095] = 16'h7817;
mem_array[22094] = 16'h3f19;
mem_array[22097] = 16'he94b;
mem_array[22096] = 16'hbe98;
mem_array[22099] = 16'h604f;
mem_array[22098] = 16'h3ebf;
mem_array[22101] = 16'h50e0;
mem_array[22100] = 16'hbdbe;
mem_array[22103] = 16'hc202;
mem_array[22102] = 16'hbd3e;
mem_array[22105] = 16'ha5bc;
mem_array[22104] = 16'hbe8f;
mem_array[22107] = 16'hb051;
mem_array[22106] = 16'hbfa5;
mem_array[22109] = 16'hdbd0;
mem_array[22108] = 16'hbf80;
mem_array[22111] = 16'h256a;
mem_array[22110] = 16'hbd32;
mem_array[22113] = 16'h20b7;
mem_array[22112] = 16'h3e18;
mem_array[22115] = 16'hcea7;
mem_array[22114] = 16'h3d2d;
mem_array[22117] = 16'h54f1;
mem_array[22116] = 16'h3ed0;
mem_array[22119] = 16'h6141;
mem_array[22118] = 16'hbe84;
mem_array[22121] = 16'h001d;
mem_array[22120] = 16'hbf97;
mem_array[22123] = 16'h6d5d;
mem_array[22122] = 16'h3e23;
mem_array[22125] = 16'ha43d;
mem_array[22124] = 16'hbefc;
mem_array[22127] = 16'h76e9;
mem_array[22126] = 16'h3f03;
mem_array[22129] = 16'h257b;
mem_array[22128] = 16'hc007;
mem_array[22131] = 16'hfe6b;
mem_array[22130] = 16'hbea4;
mem_array[22133] = 16'h85b0;
mem_array[22132] = 16'hbf11;
mem_array[22135] = 16'h3bd3;
mem_array[22134] = 16'hbf94;
mem_array[22137] = 16'hb304;
mem_array[22136] = 16'hbf08;
mem_array[22139] = 16'heab2;
mem_array[22138] = 16'hbdc4;
mem_array[22141] = 16'hffbb;
mem_array[22140] = 16'hbfad;
mem_array[22143] = 16'h4ca1;
mem_array[22142] = 16'hbd3e;
mem_array[22145] = 16'h9c7b;
mem_array[22144] = 16'h3e96;
mem_array[22147] = 16'h52d5;
mem_array[22146] = 16'hbdcb;
mem_array[22149] = 16'hd1c3;
mem_array[22148] = 16'hbebb;
mem_array[22151] = 16'h9881;
mem_array[22150] = 16'h3dc5;
mem_array[22153] = 16'h3194;
mem_array[22152] = 16'hbd91;
mem_array[22155] = 16'hd629;
mem_array[22154] = 16'h3ef0;
mem_array[22157] = 16'h4d19;
mem_array[22156] = 16'h3ee5;
mem_array[22159] = 16'h3461;
mem_array[22158] = 16'hbeb5;
mem_array[22161] = 16'hb60e;
mem_array[22160] = 16'hbd17;
mem_array[22163] = 16'h5fcb;
mem_array[22162] = 16'hbda3;
mem_array[22165] = 16'h7ca7;
mem_array[22164] = 16'hbe1c;
mem_array[22167] = 16'h76b4;
mem_array[22166] = 16'hbf98;
mem_array[22169] = 16'ha357;
mem_array[22168] = 16'hbf28;
mem_array[22171] = 16'h08a4;
mem_array[22170] = 16'hbe01;
mem_array[22173] = 16'h7450;
mem_array[22172] = 16'hbebb;
mem_array[22175] = 16'hb481;
mem_array[22174] = 16'h3d98;
mem_array[22177] = 16'h84fd;
mem_array[22176] = 16'h3e0b;
mem_array[22179] = 16'h8028;
mem_array[22178] = 16'hbcf3;
mem_array[22181] = 16'h2dc7;
mem_array[22180] = 16'hbf19;
mem_array[22183] = 16'ha02f;
mem_array[22182] = 16'h3d90;
mem_array[22185] = 16'hbdc9;
mem_array[22184] = 16'hbef1;
mem_array[22187] = 16'hdf24;
mem_array[22186] = 16'h3e49;
mem_array[22189] = 16'h7547;
mem_array[22188] = 16'hc011;
mem_array[22191] = 16'he78c;
mem_array[22190] = 16'h3d83;
mem_array[22193] = 16'h5fb4;
mem_array[22192] = 16'h3dbf;
mem_array[22195] = 16'h3722;
mem_array[22194] = 16'h3e29;
mem_array[22197] = 16'h2c54;
mem_array[22196] = 16'hbeaa;
mem_array[22199] = 16'h7d8c;
mem_array[22198] = 16'h3e65;
mem_array[22201] = 16'h7783;
mem_array[22200] = 16'hbfcf;
mem_array[22203] = 16'hd581;
mem_array[22202] = 16'h3c24;
mem_array[22205] = 16'ha166;
mem_array[22204] = 16'h3e29;
mem_array[22207] = 16'h3e3a;
mem_array[22206] = 16'h3ec3;
mem_array[22209] = 16'h9759;
mem_array[22208] = 16'hbda1;
mem_array[22211] = 16'h12d9;
mem_array[22210] = 16'hbd4a;
mem_array[22213] = 16'h4880;
mem_array[22212] = 16'h3e75;
mem_array[22215] = 16'h5824;
mem_array[22214] = 16'h3d10;
mem_array[22217] = 16'h9915;
mem_array[22216] = 16'hbee4;
mem_array[22219] = 16'h17dd;
mem_array[22218] = 16'h3eaf;
mem_array[22221] = 16'ha63c;
mem_array[22220] = 16'hbd24;
mem_array[22223] = 16'ha092;
mem_array[22222] = 16'hbd83;
mem_array[22225] = 16'h2802;
mem_array[22224] = 16'h3dbc;
mem_array[22227] = 16'hee42;
mem_array[22226] = 16'hbf7b;
mem_array[22229] = 16'h97cc;
mem_array[22228] = 16'hbfb1;
mem_array[22231] = 16'h2a10;
mem_array[22230] = 16'hbef8;
mem_array[22233] = 16'h56d1;
mem_array[22232] = 16'hbf95;
mem_array[22235] = 16'h362c;
mem_array[22234] = 16'hbdba;
mem_array[22237] = 16'h2dfc;
mem_array[22236] = 16'h3db4;
mem_array[22239] = 16'h46af;
mem_array[22238] = 16'hbcb1;
mem_array[22241] = 16'h5110;
mem_array[22240] = 16'h3e69;
mem_array[22243] = 16'h5d02;
mem_array[22242] = 16'hbd11;
mem_array[22245] = 16'h00ce;
mem_array[22244] = 16'hbe7f;
mem_array[22247] = 16'h9ba2;
mem_array[22246] = 16'h3c29;
mem_array[22249] = 16'h9545;
mem_array[22248] = 16'hc018;
mem_array[22251] = 16'he855;
mem_array[22250] = 16'hbd58;
mem_array[22253] = 16'hedcf;
mem_array[22252] = 16'hbe75;
mem_array[22255] = 16'h5f08;
mem_array[22254] = 16'h3ecd;
mem_array[22257] = 16'h65a8;
mem_array[22256] = 16'h3f0e;
mem_array[22259] = 16'hfee5;
mem_array[22258] = 16'h3e88;
mem_array[22261] = 16'h151f;
mem_array[22260] = 16'hbeed;
mem_array[22263] = 16'h0719;
mem_array[22262] = 16'h3d76;
mem_array[22265] = 16'h6c20;
mem_array[22264] = 16'h3d35;
mem_array[22267] = 16'h6d43;
mem_array[22266] = 16'h3e87;
mem_array[22269] = 16'h91ef;
mem_array[22268] = 16'h3df3;
mem_array[22271] = 16'h80ea;
mem_array[22270] = 16'h3e65;
mem_array[22273] = 16'h7f8c;
mem_array[22272] = 16'h3ea9;
mem_array[22275] = 16'hf788;
mem_array[22274] = 16'hbea9;
mem_array[22277] = 16'hefec;
mem_array[22276] = 16'hbf33;
mem_array[22279] = 16'he86f;
mem_array[22278] = 16'h3f0c;
mem_array[22281] = 16'hf5af;
mem_array[22280] = 16'hbdc4;
mem_array[22283] = 16'h0e6b;
mem_array[22282] = 16'h3cb5;
mem_array[22285] = 16'hba8f;
mem_array[22284] = 16'h3e59;
mem_array[22287] = 16'h9751;
mem_array[22286] = 16'hbf3e;
mem_array[22289] = 16'h0cba;
mem_array[22288] = 16'hbfb4;
mem_array[22291] = 16'h0d68;
mem_array[22290] = 16'hbe57;
mem_array[22293] = 16'h114c;
mem_array[22292] = 16'hbf51;
mem_array[22295] = 16'hbe59;
mem_array[22294] = 16'hbda4;
mem_array[22297] = 16'h3d65;
mem_array[22296] = 16'h3e3b;
mem_array[22299] = 16'hff81;
mem_array[22298] = 16'h3ca7;
mem_array[22301] = 16'h3b10;
mem_array[22300] = 16'hbd36;
mem_array[22303] = 16'h20d0;
mem_array[22302] = 16'h3d51;
mem_array[22305] = 16'h83ea;
mem_array[22304] = 16'hbe7b;
mem_array[22307] = 16'haa2f;
mem_array[22306] = 16'hbbf8;
mem_array[22309] = 16'h46a1;
mem_array[22308] = 16'hc035;
mem_array[22311] = 16'hf06f;
mem_array[22310] = 16'h3ecb;
mem_array[22313] = 16'habbc;
mem_array[22312] = 16'hbdbc;
mem_array[22315] = 16'h369a;
mem_array[22314] = 16'h3de9;
mem_array[22317] = 16'hd9bf;
mem_array[22316] = 16'h3efe;
mem_array[22319] = 16'he006;
mem_array[22318] = 16'hbec1;
mem_array[22321] = 16'hb689;
mem_array[22320] = 16'hbe9f;
mem_array[22323] = 16'he22e;
mem_array[22322] = 16'h3e07;
mem_array[22325] = 16'hd83b;
mem_array[22324] = 16'h3dca;
mem_array[22327] = 16'h0e4e;
mem_array[22326] = 16'h3ddd;
mem_array[22329] = 16'h8ded;
mem_array[22328] = 16'hbe0e;
mem_array[22331] = 16'h3a61;
mem_array[22330] = 16'h3d0e;
mem_array[22333] = 16'h5984;
mem_array[22332] = 16'h3edb;
mem_array[22335] = 16'h4078;
mem_array[22334] = 16'h3c48;
mem_array[22337] = 16'h3d39;
mem_array[22336] = 16'hbf8c;
mem_array[22339] = 16'hcaa7;
mem_array[22338] = 16'h3cd7;
mem_array[22341] = 16'h9780;
mem_array[22340] = 16'hbd15;
mem_array[22343] = 16'h5165;
mem_array[22342] = 16'h3cb2;
mem_array[22345] = 16'heb1f;
mem_array[22344] = 16'h3e22;
mem_array[22347] = 16'h69d5;
mem_array[22346] = 16'hbe77;
mem_array[22349] = 16'h955b;
mem_array[22348] = 16'hbfb4;
mem_array[22351] = 16'h5450;
mem_array[22350] = 16'hbe83;
mem_array[22353] = 16'h3496;
mem_array[22352] = 16'hbf90;
mem_array[22355] = 16'h289e;
mem_array[22354] = 16'h3e27;
mem_array[22357] = 16'h4432;
mem_array[22356] = 16'h3deb;
mem_array[22359] = 16'h8028;
mem_array[22358] = 16'h3e51;
mem_array[22361] = 16'h9f14;
mem_array[22360] = 16'hbd74;
mem_array[22363] = 16'ha646;
mem_array[22362] = 16'hbdac;
mem_array[22365] = 16'hf92b;
mem_array[22364] = 16'hbd44;
mem_array[22367] = 16'h9b3e;
mem_array[22366] = 16'h3e3b;
mem_array[22369] = 16'h2d69;
mem_array[22368] = 16'hbf82;
mem_array[22371] = 16'hf1ed;
mem_array[22370] = 16'h3f35;
mem_array[22373] = 16'h8cd2;
mem_array[22372] = 16'hbd89;
mem_array[22375] = 16'hc489;
mem_array[22374] = 16'h3e49;
mem_array[22377] = 16'h2cc4;
mem_array[22376] = 16'h3e1f;
mem_array[22379] = 16'h9733;
mem_array[22378] = 16'h3ed4;
mem_array[22381] = 16'h571a;
mem_array[22380] = 16'hbf4f;
mem_array[22383] = 16'h9071;
mem_array[22382] = 16'hbda1;
mem_array[22385] = 16'h5b2c;
mem_array[22384] = 16'h3e31;
mem_array[22387] = 16'h36c1;
mem_array[22386] = 16'h3e23;
mem_array[22389] = 16'h88b7;
mem_array[22388] = 16'h3d62;
mem_array[22391] = 16'h8aa4;
mem_array[22390] = 16'h3c9a;
mem_array[22393] = 16'h3278;
mem_array[22392] = 16'h3eef;
mem_array[22395] = 16'h2fff;
mem_array[22394] = 16'h3dc6;
mem_array[22397] = 16'ha84c;
mem_array[22396] = 16'hbf46;
mem_array[22399] = 16'hf07f;
mem_array[22398] = 16'h3e25;
mem_array[22401] = 16'h4a53;
mem_array[22400] = 16'h3c1f;
mem_array[22403] = 16'h6715;
mem_array[22402] = 16'hbcbd;
mem_array[22405] = 16'hb062;
mem_array[22404] = 16'hbde1;
mem_array[22407] = 16'h44d4;
mem_array[22406] = 16'h3d37;
mem_array[22409] = 16'h4d23;
mem_array[22408] = 16'hbf99;
mem_array[22411] = 16'h06d1;
mem_array[22410] = 16'hbed6;
mem_array[22413] = 16'h448d;
mem_array[22412] = 16'hbf2f;
mem_array[22415] = 16'h1a84;
mem_array[22414] = 16'h3de5;
mem_array[22417] = 16'hf984;
mem_array[22416] = 16'h3c88;
mem_array[22419] = 16'h2fd3;
mem_array[22418] = 16'hba2a;
mem_array[22421] = 16'h6e5e;
mem_array[22420] = 16'h3e12;
mem_array[22423] = 16'ha20b;
mem_array[22422] = 16'hbe38;
mem_array[22425] = 16'he3fb;
mem_array[22424] = 16'hbdd9;
mem_array[22427] = 16'hca67;
mem_array[22426] = 16'hbdec;
mem_array[22429] = 16'hc927;
mem_array[22428] = 16'hbc59;
mem_array[22431] = 16'hbe3b;
mem_array[22430] = 16'h3db6;
mem_array[22433] = 16'hb8ce;
mem_array[22432] = 16'h3e3d;
mem_array[22435] = 16'h0ee7;
mem_array[22434] = 16'h3c62;
mem_array[22437] = 16'h76c4;
mem_array[22436] = 16'h3ecc;
mem_array[22439] = 16'hf03c;
mem_array[22438] = 16'h3c92;
mem_array[22441] = 16'hfb75;
mem_array[22440] = 16'hbf37;
mem_array[22443] = 16'hc5c1;
mem_array[22442] = 16'h3e47;
mem_array[22445] = 16'he0ad;
mem_array[22444] = 16'hbf7b;
mem_array[22447] = 16'h22d3;
mem_array[22446] = 16'h3ef2;
mem_array[22449] = 16'h91bd;
mem_array[22448] = 16'hbe82;
mem_array[22451] = 16'hbe8b;
mem_array[22450] = 16'h3e06;
mem_array[22453] = 16'h40fd;
mem_array[22452] = 16'h3c84;
mem_array[22455] = 16'h8fe4;
mem_array[22454] = 16'hbd96;
mem_array[22457] = 16'h6223;
mem_array[22456] = 16'hbf54;
mem_array[22459] = 16'h7a07;
mem_array[22458] = 16'hbe50;
mem_array[22461] = 16'hde9a;
mem_array[22460] = 16'hbd92;
mem_array[22463] = 16'hf905;
mem_array[22462] = 16'h3d05;
mem_array[22465] = 16'h8db7;
mem_array[22464] = 16'h3d5c;
mem_array[22467] = 16'h4c7f;
mem_array[22466] = 16'hbe69;
mem_array[22469] = 16'h7a18;
mem_array[22468] = 16'hbfd3;
mem_array[22471] = 16'h117e;
mem_array[22470] = 16'hbe83;
mem_array[22473] = 16'hc85d;
mem_array[22472] = 16'hbe6b;
mem_array[22475] = 16'h0d03;
mem_array[22474] = 16'h3ee3;
mem_array[22477] = 16'hdb52;
mem_array[22476] = 16'h3b69;
mem_array[22479] = 16'h2c81;
mem_array[22478] = 16'hbd1b;
mem_array[22481] = 16'h691a;
mem_array[22480] = 16'h3eec;
mem_array[22483] = 16'haa08;
mem_array[22482] = 16'hbc05;
mem_array[22485] = 16'he478;
mem_array[22484] = 16'hbd08;
mem_array[22487] = 16'he26c;
mem_array[22486] = 16'hbe2a;
mem_array[22489] = 16'h74e5;
mem_array[22488] = 16'h3e28;
mem_array[22491] = 16'h11bd;
mem_array[22490] = 16'h3ed9;
mem_array[22493] = 16'h13e2;
mem_array[22492] = 16'hbe15;
mem_array[22495] = 16'ha06d;
mem_array[22494] = 16'h3e94;
mem_array[22497] = 16'h4590;
mem_array[22496] = 16'h3e27;
mem_array[22499] = 16'hf24d;
mem_array[22498] = 16'h3ebe;
mem_array[22501] = 16'h8c62;
mem_array[22500] = 16'hbdfb;
mem_array[22503] = 16'hba4f;
mem_array[22502] = 16'h3da0;
mem_array[22505] = 16'hb9c2;
mem_array[22504] = 16'hc033;
mem_array[22507] = 16'h4534;
mem_array[22506] = 16'h3d3b;
mem_array[22509] = 16'h2c34;
mem_array[22508] = 16'h3d8d;
mem_array[22511] = 16'h59ac;
mem_array[22510] = 16'h3e84;
mem_array[22513] = 16'h97ab;
mem_array[22512] = 16'hbe18;
mem_array[22515] = 16'h555b;
mem_array[22514] = 16'hbe70;
mem_array[22517] = 16'h0902;
mem_array[22516] = 16'hbeb0;
mem_array[22519] = 16'hd430;
mem_array[22518] = 16'hbec1;
mem_array[22521] = 16'h133c;
mem_array[22520] = 16'hbcc8;
mem_array[22523] = 16'hf5fe;
mem_array[22522] = 16'hbcf9;
mem_array[22525] = 16'h4dc1;
mem_array[22524] = 16'h3d5d;
mem_array[22527] = 16'hea63;
mem_array[22526] = 16'hbdbb;
mem_array[22529] = 16'h2689;
mem_array[22528] = 16'hc010;
mem_array[22531] = 16'h01d7;
mem_array[22530] = 16'h3e20;
mem_array[22533] = 16'hf907;
mem_array[22532] = 16'hbf0b;
mem_array[22535] = 16'h34a7;
mem_array[22534] = 16'h3eb7;
mem_array[22537] = 16'h1d33;
mem_array[22536] = 16'h3de0;
mem_array[22539] = 16'h8f58;
mem_array[22538] = 16'h3e67;
mem_array[22541] = 16'hd40c;
mem_array[22540] = 16'h3e91;
mem_array[22543] = 16'h5b39;
mem_array[22542] = 16'h3e4b;
mem_array[22545] = 16'h1125;
mem_array[22544] = 16'hbe2c;
mem_array[22547] = 16'h3094;
mem_array[22546] = 16'hbda5;
mem_array[22549] = 16'h2269;
mem_array[22548] = 16'h3e31;
mem_array[22551] = 16'hdae8;
mem_array[22550] = 16'h3ef8;
mem_array[22553] = 16'h0716;
mem_array[22552] = 16'h3e8e;
mem_array[22555] = 16'h10c7;
mem_array[22554] = 16'h3e7a;
mem_array[22557] = 16'h7d96;
mem_array[22556] = 16'h3eaa;
mem_array[22559] = 16'h0705;
mem_array[22558] = 16'h3ec1;
mem_array[22561] = 16'h0194;
mem_array[22560] = 16'hbece;
mem_array[22563] = 16'hfa64;
mem_array[22562] = 16'hbeb1;
mem_array[22565] = 16'h7336;
mem_array[22564] = 16'hbf47;
mem_array[22567] = 16'haa18;
mem_array[22566] = 16'hbeed;
mem_array[22569] = 16'hb273;
mem_array[22568] = 16'hbeab;
mem_array[22571] = 16'h0b78;
mem_array[22570] = 16'h3ea0;
mem_array[22573] = 16'hd28f;
mem_array[22572] = 16'hbe25;
mem_array[22575] = 16'h25ce;
mem_array[22574] = 16'h3d3e;
mem_array[22577] = 16'h68af;
mem_array[22576] = 16'hbea1;
mem_array[22579] = 16'h6dcc;
mem_array[22578] = 16'hbe28;
mem_array[22581] = 16'hc696;
mem_array[22580] = 16'h3c78;
mem_array[22583] = 16'h1525;
mem_array[22582] = 16'h3c9a;
mem_array[22585] = 16'hcf09;
mem_array[22584] = 16'h3bd2;
mem_array[22587] = 16'hd1e7;
mem_array[22586] = 16'h3e0a;
mem_array[22589] = 16'h4bd0;
mem_array[22588] = 16'hbfe8;
mem_array[22591] = 16'h2304;
mem_array[22590] = 16'h3e80;
mem_array[22593] = 16'h8c40;
mem_array[22592] = 16'hbe88;
mem_array[22595] = 16'h0f7a;
mem_array[22594] = 16'hbd93;
mem_array[22597] = 16'h4af4;
mem_array[22596] = 16'hbe93;
mem_array[22599] = 16'h0d5b;
mem_array[22598] = 16'h3de9;
mem_array[22601] = 16'h1a04;
mem_array[22600] = 16'h3ec8;
mem_array[22603] = 16'h0efd;
mem_array[22602] = 16'h3e07;
mem_array[22605] = 16'h3e0d;
mem_array[22604] = 16'h3e43;
mem_array[22607] = 16'hdb55;
mem_array[22606] = 16'hbe80;
mem_array[22609] = 16'h7c4e;
mem_array[22608] = 16'h3ebd;
mem_array[22611] = 16'h7bbd;
mem_array[22610] = 16'hbf35;
mem_array[22613] = 16'hf064;
mem_array[22612] = 16'h3db9;
mem_array[22615] = 16'hf7c9;
mem_array[22614] = 16'h3e40;
mem_array[22617] = 16'h1393;
mem_array[22616] = 16'h3eb1;
mem_array[22619] = 16'h0201;
mem_array[22618] = 16'h3c25;
mem_array[22621] = 16'hb574;
mem_array[22620] = 16'h3e7d;
mem_array[22623] = 16'h180b;
mem_array[22622] = 16'hbf76;
mem_array[22625] = 16'he496;
mem_array[22624] = 16'h3ea3;
mem_array[22627] = 16'he037;
mem_array[22626] = 16'hbf73;
mem_array[22629] = 16'hb3ba;
mem_array[22628] = 16'hbef2;
mem_array[22631] = 16'had44;
mem_array[22630] = 16'h3df9;
mem_array[22633] = 16'h24df;
mem_array[22632] = 16'h3e22;
mem_array[22635] = 16'hba6d;
mem_array[22634] = 16'hbdbc;
mem_array[22637] = 16'he9e4;
mem_array[22636] = 16'hbe0c;
mem_array[22639] = 16'h9df5;
mem_array[22638] = 16'hbeae;
mem_array[22641] = 16'hd738;
mem_array[22640] = 16'hbcc0;
mem_array[22643] = 16'ha61b;
mem_array[22642] = 16'h3d07;
mem_array[22645] = 16'hf7ca;
mem_array[22644] = 16'h3a76;
mem_array[22647] = 16'hf3ed;
mem_array[22646] = 16'h3cec;
mem_array[22649] = 16'hdc0e;
mem_array[22648] = 16'hbfa2;
mem_array[22651] = 16'h2103;
mem_array[22650] = 16'h3d89;
mem_array[22653] = 16'hea5f;
mem_array[22652] = 16'h3c5d;
mem_array[22655] = 16'h71a2;
mem_array[22654] = 16'hbefc;
mem_array[22657] = 16'h57c6;
mem_array[22656] = 16'hbe4f;
mem_array[22659] = 16'h4968;
mem_array[22658] = 16'hbe0d;
mem_array[22661] = 16'h3019;
mem_array[22660] = 16'h3e03;
mem_array[22663] = 16'h036d;
mem_array[22662] = 16'h3e0b;
mem_array[22665] = 16'hc8a7;
mem_array[22664] = 16'h3e2b;
mem_array[22667] = 16'h24d6;
mem_array[22666] = 16'hbe50;
mem_array[22669] = 16'hbbcd;
mem_array[22668] = 16'h3ee0;
mem_array[22671] = 16'h546f;
mem_array[22670] = 16'hc001;
mem_array[22673] = 16'h2146;
mem_array[22672] = 16'hbccf;
mem_array[22675] = 16'h2641;
mem_array[22674] = 16'hbd26;
mem_array[22677] = 16'h2d1f;
mem_array[22676] = 16'h3ecb;
mem_array[22679] = 16'h8e0a;
mem_array[22678] = 16'hbe6a;
mem_array[22681] = 16'hccae;
mem_array[22680] = 16'h3e2f;
mem_array[22683] = 16'h54e8;
mem_array[22682] = 16'hbf36;
mem_array[22685] = 16'h35dd;
mem_array[22684] = 16'hbe92;
mem_array[22687] = 16'hb8a3;
mem_array[22686] = 16'hbfb6;
mem_array[22689] = 16'hf4c1;
mem_array[22688] = 16'h3cbf;
mem_array[22691] = 16'h526d;
mem_array[22690] = 16'h3db0;
mem_array[22693] = 16'h3ecd;
mem_array[22692] = 16'h3ea6;
mem_array[22695] = 16'hdc2a;
mem_array[22694] = 16'h3e37;
mem_array[22697] = 16'h2711;
mem_array[22696] = 16'hbd6a;
mem_array[22699] = 16'hbb71;
mem_array[22698] = 16'h3dc9;
mem_array[22701] = 16'h64dd;
mem_array[22700] = 16'hbd88;
mem_array[22703] = 16'h0e3d;
mem_array[22702] = 16'h3cd2;
mem_array[22705] = 16'h4cd9;
mem_array[22704] = 16'hbe3f;
mem_array[22707] = 16'h50f6;
mem_array[22706] = 16'hbf11;
mem_array[22709] = 16'hb89c;
mem_array[22708] = 16'hbf76;
mem_array[22711] = 16'h971f;
mem_array[22710] = 16'h3e6d;
mem_array[22713] = 16'h360d;
mem_array[22712] = 16'hbe06;
mem_array[22715] = 16'h9718;
mem_array[22714] = 16'hbe99;
mem_array[22717] = 16'h2879;
mem_array[22716] = 16'hbd4b;
mem_array[22719] = 16'h991b;
mem_array[22718] = 16'hbec5;
mem_array[22721] = 16'hcf72;
mem_array[22720] = 16'hbcc6;
mem_array[22723] = 16'ha05a;
mem_array[22722] = 16'h3d6f;
mem_array[22725] = 16'he979;
mem_array[22724] = 16'hbe18;
mem_array[22727] = 16'hba2c;
mem_array[22726] = 16'hbe2d;
mem_array[22729] = 16'hf8a6;
mem_array[22728] = 16'h3d5f;
mem_array[22731] = 16'h6c9d;
mem_array[22730] = 16'hbea0;
mem_array[22733] = 16'h7aa5;
mem_array[22732] = 16'h3da8;
mem_array[22735] = 16'h03e9;
mem_array[22734] = 16'h3d1a;
mem_array[22737] = 16'h45dc;
mem_array[22736] = 16'h3e36;
mem_array[22739] = 16'hf62e;
mem_array[22738] = 16'hbee7;
mem_array[22741] = 16'h1a1b;
mem_array[22740] = 16'h3e28;
mem_array[22743] = 16'h12c0;
mem_array[22742] = 16'hbf1e;
mem_array[22745] = 16'hfdaa;
mem_array[22744] = 16'hbe00;
mem_array[22747] = 16'ha4dd;
mem_array[22746] = 16'hbfa8;
mem_array[22749] = 16'hbd09;
mem_array[22748] = 16'hbc95;
mem_array[22751] = 16'h6b8b;
mem_array[22750] = 16'h3d88;
mem_array[22753] = 16'h1005;
mem_array[22752] = 16'hbd7c;
mem_array[22755] = 16'hddf9;
mem_array[22754] = 16'h3e50;
mem_array[22757] = 16'ha619;
mem_array[22756] = 16'hbbc1;
mem_array[22759] = 16'h1734;
mem_array[22758] = 16'hbdb6;
mem_array[22761] = 16'h50a5;
mem_array[22760] = 16'h3cb1;
mem_array[22763] = 16'h7ecc;
mem_array[22762] = 16'hbcfb;
mem_array[22765] = 16'h30c6;
mem_array[22764] = 16'hbe08;
mem_array[22767] = 16'h3b4e;
mem_array[22766] = 16'hbf01;
mem_array[22769] = 16'hdc67;
mem_array[22768] = 16'hbec0;
mem_array[22771] = 16'h6d7e;
mem_array[22770] = 16'h3e80;
mem_array[22773] = 16'h9561;
mem_array[22772] = 16'hbdd4;
mem_array[22775] = 16'hc459;
mem_array[22774] = 16'hbd62;
mem_array[22777] = 16'h473e;
mem_array[22776] = 16'h3e9c;
mem_array[22779] = 16'h1ae1;
mem_array[22778] = 16'hbf45;
mem_array[22781] = 16'h723f;
mem_array[22780] = 16'h3e29;
mem_array[22783] = 16'hc017;
mem_array[22782] = 16'h3cdf;
mem_array[22785] = 16'h71df;
mem_array[22784] = 16'hbd84;
mem_array[22787] = 16'heba0;
mem_array[22786] = 16'hbe26;
mem_array[22789] = 16'he7a8;
mem_array[22788] = 16'hbe28;
mem_array[22791] = 16'h1b6a;
mem_array[22790] = 16'h3dad;
mem_array[22793] = 16'h6e7f;
mem_array[22792] = 16'hbe01;
mem_array[22795] = 16'hc97a;
mem_array[22794] = 16'hbeac;
mem_array[22797] = 16'h8f8c;
mem_array[22796] = 16'hbdba;
mem_array[22799] = 16'h8894;
mem_array[22798] = 16'hbe30;
mem_array[22801] = 16'h3895;
mem_array[22800] = 16'h3dc3;
mem_array[22803] = 16'h9f62;
mem_array[22802] = 16'hbdb1;
mem_array[22805] = 16'h19d4;
mem_array[22804] = 16'hbe19;
mem_array[22807] = 16'h879e;
mem_array[22806] = 16'hbfa7;
mem_array[22809] = 16'h2b93;
mem_array[22808] = 16'h3e10;
mem_array[22811] = 16'hf4df;
mem_array[22810] = 16'hbe61;
mem_array[22813] = 16'h7fce;
mem_array[22812] = 16'h3d56;
mem_array[22815] = 16'h7784;
mem_array[22814] = 16'h3e80;
mem_array[22817] = 16'h9257;
mem_array[22816] = 16'hbec6;
mem_array[22819] = 16'hac1b;
mem_array[22818] = 16'hbd16;
mem_array[22821] = 16'hd0cd;
mem_array[22820] = 16'hbdf5;
mem_array[22823] = 16'h99f7;
mem_array[22822] = 16'h3c3e;
mem_array[22825] = 16'he9b7;
mem_array[22824] = 16'hbc64;
mem_array[22827] = 16'h56c9;
mem_array[22826] = 16'hbe2c;
mem_array[22829] = 16'h5d37;
mem_array[22828] = 16'hbedf;
mem_array[22831] = 16'ha2f8;
mem_array[22830] = 16'h3da7;
mem_array[22833] = 16'hf293;
mem_array[22832] = 16'h3d3d;
mem_array[22835] = 16'h53e6;
mem_array[22834] = 16'hbcb1;
mem_array[22837] = 16'he980;
mem_array[22836] = 16'h3eb3;
mem_array[22839] = 16'h4424;
mem_array[22838] = 16'hbe50;
mem_array[22841] = 16'h175b;
mem_array[22840] = 16'h3e99;
mem_array[22843] = 16'h2943;
mem_array[22842] = 16'h3d07;
mem_array[22845] = 16'h0ba2;
mem_array[22844] = 16'h3d43;
mem_array[22847] = 16'h9f0f;
mem_array[22846] = 16'hbd76;
mem_array[22849] = 16'h3358;
mem_array[22848] = 16'h3e11;
mem_array[22851] = 16'hfea5;
mem_array[22850] = 16'h3dea;
mem_array[22853] = 16'h47cc;
mem_array[22852] = 16'hbdec;
mem_array[22855] = 16'hd3ab;
mem_array[22854] = 16'hbefc;
mem_array[22857] = 16'hc60e;
mem_array[22856] = 16'h3e15;
mem_array[22859] = 16'h9589;
mem_array[22858] = 16'hbd72;
mem_array[22861] = 16'hb2e4;
mem_array[22860] = 16'h3d36;
mem_array[22863] = 16'h30ec;
mem_array[22862] = 16'h3da8;
mem_array[22865] = 16'h1c7f;
mem_array[22864] = 16'h3d13;
mem_array[22867] = 16'hf957;
mem_array[22866] = 16'hbea9;
mem_array[22869] = 16'h7716;
mem_array[22868] = 16'hbcca;
mem_array[22871] = 16'hc3dc;
mem_array[22870] = 16'hbd4f;
mem_array[22873] = 16'h4689;
mem_array[22872] = 16'hbc1a;
mem_array[22875] = 16'h30f1;
mem_array[22874] = 16'hbd55;
mem_array[22877] = 16'h90d8;
mem_array[22876] = 16'hbd35;
mem_array[22879] = 16'h8fd3;
mem_array[22878] = 16'hbec9;
mem_array[22881] = 16'hc08d;
mem_array[22880] = 16'hbd79;
mem_array[22883] = 16'h9e7f;
mem_array[22882] = 16'h3d0a;
mem_array[22885] = 16'hcd55;
mem_array[22884] = 16'hbc6f;
mem_array[22887] = 16'h0c45;
mem_array[22886] = 16'hbea8;
mem_array[22889] = 16'hd95b;
mem_array[22888] = 16'hbeb5;
mem_array[22891] = 16'hb96c;
mem_array[22890] = 16'h3ddb;
mem_array[22893] = 16'h479a;
mem_array[22892] = 16'h3e78;
mem_array[22895] = 16'h05ad;
mem_array[22894] = 16'h3d8f;
mem_array[22897] = 16'he5be;
mem_array[22896] = 16'h3ed9;
mem_array[22899] = 16'hf9ee;
mem_array[22898] = 16'h3eba;
mem_array[22901] = 16'h7d25;
mem_array[22900] = 16'h3da1;
mem_array[22903] = 16'hc8d2;
mem_array[22902] = 16'h3cb5;
mem_array[22905] = 16'hc025;
mem_array[22904] = 16'h3e34;
mem_array[22907] = 16'he26f;
mem_array[22906] = 16'hbe44;
mem_array[22909] = 16'h59c3;
mem_array[22908] = 16'h3e24;
mem_array[22911] = 16'hdacc;
mem_array[22910] = 16'hbe6c;
mem_array[22913] = 16'hf11c;
mem_array[22912] = 16'hbe3c;
mem_array[22915] = 16'hee22;
mem_array[22914] = 16'hbf2b;
mem_array[22917] = 16'hb360;
mem_array[22916] = 16'hbe08;
mem_array[22919] = 16'habd6;
mem_array[22918] = 16'h3e94;
mem_array[22921] = 16'hda74;
mem_array[22920] = 16'hbedb;
mem_array[22923] = 16'h01ba;
mem_array[22922] = 16'hbdae;
mem_array[22925] = 16'h7c38;
mem_array[22924] = 16'hbd4d;
mem_array[22927] = 16'he525;
mem_array[22926] = 16'hbe1e;
mem_array[22929] = 16'h8166;
mem_array[22928] = 16'hbe4e;
mem_array[22931] = 16'h6172;
mem_array[22930] = 16'hbd8d;
mem_array[22933] = 16'h1440;
mem_array[22932] = 16'hbe2e;
mem_array[22935] = 16'h2fab;
mem_array[22934] = 16'hbce7;
mem_array[22937] = 16'hc2db;
mem_array[22936] = 16'hbd84;
mem_array[22939] = 16'h52d1;
mem_array[22938] = 16'hbf75;
mem_array[22941] = 16'hd8dd;
mem_array[22940] = 16'hbe0c;
mem_array[22943] = 16'h4aa0;
mem_array[22942] = 16'hbd0c;
mem_array[22945] = 16'hfe21;
mem_array[22944] = 16'hbcf6;
mem_array[22947] = 16'h8bed;
mem_array[22946] = 16'hbc75;
mem_array[22949] = 16'h5ebd;
mem_array[22948] = 16'hbec0;
mem_array[22951] = 16'hc3ec;
mem_array[22950] = 16'h3de2;
mem_array[22953] = 16'haf76;
mem_array[22952] = 16'h3e90;
mem_array[22955] = 16'h3f71;
mem_array[22954] = 16'h3d9b;
mem_array[22957] = 16'h0fad;
mem_array[22956] = 16'h3e4a;
mem_array[22959] = 16'h8a3d;
mem_array[22958] = 16'h3e26;
mem_array[22961] = 16'hb0d7;
mem_array[22960] = 16'h3caa;
mem_array[22963] = 16'hc2a8;
mem_array[22962] = 16'h3e14;
mem_array[22965] = 16'h87b1;
mem_array[22964] = 16'h3e4d;
mem_array[22967] = 16'h7723;
mem_array[22966] = 16'h3dcf;
mem_array[22969] = 16'h85c6;
mem_array[22968] = 16'h3d66;
mem_array[22971] = 16'h39f9;
mem_array[22970] = 16'hbe78;
mem_array[22973] = 16'h93fe;
mem_array[22972] = 16'hbced;
mem_array[22975] = 16'ha579;
mem_array[22974] = 16'hbfa6;
mem_array[22977] = 16'h71ae;
mem_array[22976] = 16'hbd78;
mem_array[22979] = 16'h6764;
mem_array[22978] = 16'hbdb4;
mem_array[22981] = 16'h0128;
mem_array[22980] = 16'hbe88;
mem_array[22983] = 16'h62ad;
mem_array[22982] = 16'hbecb;
mem_array[22985] = 16'he7f6;
mem_array[22984] = 16'hbe2d;
mem_array[22987] = 16'h18e1;
mem_array[22986] = 16'hbe73;
mem_array[22989] = 16'h0a57;
mem_array[22988] = 16'h3e4b;
mem_array[22991] = 16'he627;
mem_array[22990] = 16'hbee5;
mem_array[22993] = 16'h0c75;
mem_array[22992] = 16'hbf07;
mem_array[22995] = 16'h4737;
mem_array[22994] = 16'hbdb8;
mem_array[22997] = 16'hd2e8;
mem_array[22996] = 16'h3c68;
mem_array[22999] = 16'h1ec7;
mem_array[22998] = 16'hbd14;
mem_array[23001] = 16'h0b45;
mem_array[23000] = 16'h3c72;
mem_array[23003] = 16'hb896;
mem_array[23002] = 16'hbd8a;
mem_array[23005] = 16'hefef;
mem_array[23004] = 16'h3e0a;
mem_array[23007] = 16'h17e2;
mem_array[23006] = 16'h3da4;
mem_array[23009] = 16'h1fbe;
mem_array[23008] = 16'hbcb4;
mem_array[23011] = 16'hd3ec;
mem_array[23010] = 16'h3d48;
mem_array[23013] = 16'he844;
mem_array[23012] = 16'h3e28;
mem_array[23015] = 16'h117d;
mem_array[23014] = 16'h3d0f;
mem_array[23017] = 16'h99b2;
mem_array[23016] = 16'hbe24;
mem_array[23019] = 16'ha05c;
mem_array[23018] = 16'hbe0d;
mem_array[23021] = 16'hd6d2;
mem_array[23020] = 16'h3d5b;
mem_array[23023] = 16'hcc6f;
mem_array[23022] = 16'h3df0;
mem_array[23025] = 16'h0dbf;
mem_array[23024] = 16'h3e13;
mem_array[23027] = 16'he1ba;
mem_array[23026] = 16'hbdb8;
mem_array[23029] = 16'hb7d8;
mem_array[23028] = 16'hbf0f;
mem_array[23031] = 16'h67b8;
mem_array[23030] = 16'hbf23;
mem_array[23033] = 16'hb438;
mem_array[23032] = 16'hbbe5;
mem_array[23035] = 16'h396e;
mem_array[23034] = 16'hbfdc;
mem_array[23037] = 16'hc5c4;
mem_array[23036] = 16'hbe9a;
mem_array[23039] = 16'hffc7;
mem_array[23038] = 16'hbe47;
mem_array[23041] = 16'h39aa;
mem_array[23040] = 16'hbeb7;
mem_array[23043] = 16'hc2b6;
mem_array[23042] = 16'hbd7a;
mem_array[23045] = 16'ha96d;
mem_array[23044] = 16'hbe73;
mem_array[23047] = 16'h9258;
mem_array[23046] = 16'hbe89;
mem_array[23049] = 16'h0449;
mem_array[23048] = 16'h3e47;
mem_array[23051] = 16'h5ee8;
mem_array[23050] = 16'hbe4a;
mem_array[23053] = 16'h27b1;
mem_array[23052] = 16'hbe3d;
mem_array[23055] = 16'h3f58;
mem_array[23054] = 16'hbe18;
mem_array[23057] = 16'h16a2;
mem_array[23056] = 16'h3d25;
mem_array[23059] = 16'h40ff;
mem_array[23058] = 16'h3e61;
mem_array[23061] = 16'h001f;
mem_array[23060] = 16'h3c04;
mem_array[23063] = 16'he6d4;
mem_array[23062] = 16'h3d50;
mem_array[23065] = 16'h022d;
mem_array[23064] = 16'h3c01;
mem_array[23067] = 16'ha061;
mem_array[23066] = 16'hbe68;
mem_array[23069] = 16'h95c8;
mem_array[23068] = 16'hbe7f;
mem_array[23071] = 16'h8f73;
mem_array[23070] = 16'h3dc4;
mem_array[23073] = 16'h462a;
mem_array[23072] = 16'hbf84;
mem_array[23075] = 16'hfcf3;
mem_array[23074] = 16'h3d99;
mem_array[23077] = 16'hd39e;
mem_array[23076] = 16'hbc95;
mem_array[23079] = 16'h351a;
mem_array[23078] = 16'hbe44;
mem_array[23081] = 16'he969;
mem_array[23080] = 16'h3f26;
mem_array[23083] = 16'hd942;
mem_array[23082] = 16'h3e57;
mem_array[23085] = 16'hd777;
mem_array[23084] = 16'hbcc9;
mem_array[23087] = 16'h8ac5;
mem_array[23086] = 16'hbd58;
mem_array[23089] = 16'h544e;
mem_array[23088] = 16'hbebe;
mem_array[23091] = 16'h2c2c;
mem_array[23090] = 16'hbebf;
mem_array[23093] = 16'had36;
mem_array[23092] = 16'h3dc5;
mem_array[23095] = 16'hb338;
mem_array[23094] = 16'hc006;
mem_array[23097] = 16'h6a02;
mem_array[23096] = 16'hbe5f;
mem_array[23099] = 16'hac82;
mem_array[23098] = 16'hbe3d;
mem_array[23101] = 16'h881e;
mem_array[23100] = 16'h3f24;
mem_array[23103] = 16'h28f7;
mem_array[23102] = 16'h3e50;
mem_array[23105] = 16'hae3c;
mem_array[23104] = 16'hbd18;
mem_array[23107] = 16'hf49a;
mem_array[23106] = 16'h3dd2;
mem_array[23109] = 16'h5a15;
mem_array[23108] = 16'h3d1d;
mem_array[23111] = 16'h745f;
mem_array[23110] = 16'hbe4b;
mem_array[23113] = 16'hee5f;
mem_array[23112] = 16'hbe05;
mem_array[23115] = 16'hbd73;
mem_array[23114] = 16'hbe47;
mem_array[23117] = 16'ha7cb;
mem_array[23116] = 16'hbf12;
mem_array[23119] = 16'h2a79;
mem_array[23118] = 16'hbe6d;
mem_array[23121] = 16'hdc61;
mem_array[23120] = 16'h3d28;
mem_array[23123] = 16'hb029;
mem_array[23122] = 16'hbc56;
mem_array[23125] = 16'h7a40;
mem_array[23124] = 16'h3e96;
mem_array[23127] = 16'hea11;
mem_array[23126] = 16'hbe62;
mem_array[23129] = 16'h354b;
mem_array[23128] = 16'hbdc9;
mem_array[23131] = 16'h1450;
mem_array[23130] = 16'h3e06;
mem_array[23133] = 16'h6d2b;
mem_array[23132] = 16'hbfb4;
mem_array[23135] = 16'hb3a0;
mem_array[23134] = 16'h3ef7;
mem_array[23137] = 16'hde8e;
mem_array[23136] = 16'h3ebd;
mem_array[23139] = 16'hf703;
mem_array[23138] = 16'h3d64;
mem_array[23141] = 16'hd21c;
mem_array[23140] = 16'h3dd1;
mem_array[23143] = 16'h659d;
mem_array[23142] = 16'h3e9c;
mem_array[23145] = 16'h0d12;
mem_array[23144] = 16'h3e77;
mem_array[23147] = 16'h89a2;
mem_array[23146] = 16'hbda4;
mem_array[23149] = 16'hfdac;
mem_array[23148] = 16'h3eb7;
mem_array[23151] = 16'hdb71;
mem_array[23150] = 16'h3d7b;
mem_array[23153] = 16'h26e7;
mem_array[23152] = 16'h3d87;
mem_array[23155] = 16'ha402;
mem_array[23154] = 16'hc037;
mem_array[23157] = 16'h7c00;
mem_array[23156] = 16'h3d84;
mem_array[23159] = 16'hd029;
mem_array[23158] = 16'hbe7d;
mem_array[23161] = 16'h5e67;
mem_array[23160] = 16'h3e64;
mem_array[23163] = 16'h1aa2;
mem_array[23162] = 16'hbeca;
mem_array[23165] = 16'h0240;
mem_array[23164] = 16'hbecc;
mem_array[23167] = 16'ha5b1;
mem_array[23166] = 16'h3e05;
mem_array[23169] = 16'h478a;
mem_array[23168] = 16'h3e6b;
mem_array[23171] = 16'h149c;
mem_array[23170] = 16'hbf00;
mem_array[23173] = 16'h90c4;
mem_array[23172] = 16'hbeee;
mem_array[23175] = 16'hdb2f;
mem_array[23174] = 16'hbeb8;
mem_array[23177] = 16'h941d;
mem_array[23176] = 16'hbf00;
mem_array[23179] = 16'hdea1;
mem_array[23178] = 16'hbf3d;
mem_array[23181] = 16'hf89c;
mem_array[23180] = 16'hbd7d;
mem_array[23183] = 16'haa9d;
mem_array[23182] = 16'hbd08;
mem_array[23185] = 16'hdbdf;
mem_array[23184] = 16'h3e66;
mem_array[23187] = 16'h6a54;
mem_array[23186] = 16'hbcc6;
mem_array[23189] = 16'hf724;
mem_array[23188] = 16'h3d1c;
mem_array[23191] = 16'h5960;
mem_array[23190] = 16'h3e51;
mem_array[23193] = 16'h1d62;
mem_array[23192] = 16'hbfab;
mem_array[23195] = 16'h305a;
mem_array[23194] = 16'h3d5b;
mem_array[23197] = 16'h71d0;
mem_array[23196] = 16'h3c15;
mem_array[23199] = 16'h6472;
mem_array[23198] = 16'hbecc;
mem_array[23201] = 16'h3921;
mem_array[23200] = 16'hbe45;
mem_array[23203] = 16'h5075;
mem_array[23202] = 16'h3ea0;
mem_array[23205] = 16'hc320;
mem_array[23204] = 16'h3d80;
mem_array[23207] = 16'hfb9f;
mem_array[23206] = 16'h3f1f;
mem_array[23209] = 16'h4ada;
mem_array[23208] = 16'hbcaa;
mem_array[23211] = 16'h3943;
mem_array[23210] = 16'hbf18;
mem_array[23213] = 16'h41a0;
mem_array[23212] = 16'hbf0e;
mem_array[23215] = 16'h3c81;
mem_array[23214] = 16'hc01b;
mem_array[23217] = 16'hbe1e;
mem_array[23216] = 16'hbcf6;
mem_array[23219] = 16'hd867;
mem_array[23218] = 16'hbd55;
mem_array[23221] = 16'haf21;
mem_array[23220] = 16'h3e39;
mem_array[23223] = 16'hfcd6;
mem_array[23222] = 16'hbf11;
mem_array[23225] = 16'h775b;
mem_array[23224] = 16'hbe79;
mem_array[23227] = 16'h7f7d;
mem_array[23226] = 16'h3eeb;
mem_array[23229] = 16'h540b;
mem_array[23228] = 16'hbe71;
mem_array[23231] = 16'hbac5;
mem_array[23230] = 16'hbf13;
mem_array[23233] = 16'hfd8b;
mem_array[23232] = 16'hbe52;
mem_array[23235] = 16'h952a;
mem_array[23234] = 16'hbf23;
mem_array[23237] = 16'hb963;
mem_array[23236] = 16'h3dab;
mem_array[23239] = 16'h4d3c;
mem_array[23238] = 16'hbf83;
mem_array[23241] = 16'h3dd6;
mem_array[23240] = 16'hbb41;
mem_array[23243] = 16'hb377;
mem_array[23242] = 16'hbdc0;
mem_array[23245] = 16'h3016;
mem_array[23244] = 16'h3f1f;
mem_array[23247] = 16'h0400;
mem_array[23246] = 16'hbe09;
mem_array[23249] = 16'hb9ab;
mem_array[23248] = 16'hbe06;
mem_array[23251] = 16'hc59b;
mem_array[23250] = 16'h3ecf;
mem_array[23253] = 16'hf1f0;
mem_array[23252] = 16'hbf47;
mem_array[23255] = 16'hf95a;
mem_array[23254] = 16'hbe2f;
mem_array[23257] = 16'h67f6;
mem_array[23256] = 16'hbf30;
mem_array[23259] = 16'hdbc6;
mem_array[23258] = 16'hbf5f;
mem_array[23261] = 16'hc38b;
mem_array[23260] = 16'hbb39;
mem_array[23263] = 16'h8672;
mem_array[23262] = 16'h3d77;
mem_array[23265] = 16'h8360;
mem_array[23264] = 16'hbf40;
mem_array[23267] = 16'h7be4;
mem_array[23266] = 16'h3f35;
mem_array[23269] = 16'h3d8f;
mem_array[23268] = 16'h3e5c;
mem_array[23271] = 16'h431c;
mem_array[23270] = 16'hbf2a;
mem_array[23273] = 16'h3ee6;
mem_array[23272] = 16'hbeda;
mem_array[23275] = 16'hcfe6;
mem_array[23274] = 16'hc004;
mem_array[23277] = 16'h6e54;
mem_array[23276] = 16'h3ee6;
mem_array[23279] = 16'hfefe;
mem_array[23278] = 16'h3b1e;
mem_array[23281] = 16'h89bc;
mem_array[23280] = 16'h3ee7;
mem_array[23283] = 16'h161b;
mem_array[23282] = 16'hbe43;
mem_array[23285] = 16'h1d9a;
mem_array[23284] = 16'h3ddd;
mem_array[23287] = 16'hb17d;
mem_array[23286] = 16'h3ec4;
mem_array[23289] = 16'h0d73;
mem_array[23288] = 16'hbedd;
mem_array[23291] = 16'h51b9;
mem_array[23290] = 16'hbe70;
mem_array[23293] = 16'h4c5f;
mem_array[23292] = 16'h3e9e;
mem_array[23295] = 16'h12f9;
mem_array[23294] = 16'hbf53;
mem_array[23297] = 16'h23be;
mem_array[23296] = 16'h3e38;
mem_array[23299] = 16'h4b6f;
mem_array[23298] = 16'hbf5c;
mem_array[23301] = 16'h70a8;
mem_array[23300] = 16'h3d38;
mem_array[23303] = 16'h9891;
mem_array[23302] = 16'hbc10;
mem_array[23305] = 16'hc12f;
mem_array[23304] = 16'h3f1a;
mem_array[23307] = 16'h23e0;
mem_array[23306] = 16'h3f17;
mem_array[23309] = 16'h73e6;
mem_array[23308] = 16'h3f05;
mem_array[23311] = 16'hb699;
mem_array[23310] = 16'h3ead;
mem_array[23313] = 16'h1782;
mem_array[23312] = 16'hbf6e;
mem_array[23315] = 16'h596b;
mem_array[23314] = 16'h3e90;
mem_array[23317] = 16'hd169;
mem_array[23316] = 16'hbf46;
mem_array[23319] = 16'h292c;
mem_array[23318] = 16'hbe61;
mem_array[23321] = 16'h3dbe;
mem_array[23320] = 16'h3ef7;
mem_array[23323] = 16'hb09c;
mem_array[23322] = 16'h3c74;
mem_array[23325] = 16'hb01b;
mem_array[23324] = 16'hbf73;
mem_array[23327] = 16'h4851;
mem_array[23326] = 16'h3ed7;
mem_array[23329] = 16'h3598;
mem_array[23328] = 16'h3daa;
mem_array[23331] = 16'h1c92;
mem_array[23330] = 16'hbf0b;
mem_array[23333] = 16'h6554;
mem_array[23332] = 16'hbf1c;
mem_array[23335] = 16'haaa7;
mem_array[23334] = 16'hbf5c;
mem_array[23337] = 16'he15a;
mem_array[23336] = 16'h3eca;
mem_array[23339] = 16'hd7ee;
mem_array[23338] = 16'h3dad;
mem_array[23341] = 16'heee7;
mem_array[23340] = 16'h3f2b;
mem_array[23343] = 16'h5220;
mem_array[23342] = 16'h3e35;
mem_array[23345] = 16'hb888;
mem_array[23344] = 16'h3f2e;
mem_array[23347] = 16'h5d3d;
mem_array[23346] = 16'hbeb2;
mem_array[23349] = 16'h57d9;
mem_array[23348] = 16'h3f14;
mem_array[23351] = 16'h9d11;
mem_array[23350] = 16'hbed6;
mem_array[23353] = 16'h42d6;
mem_array[23352] = 16'h3f16;
mem_array[23355] = 16'hfc3e;
mem_array[23354] = 16'hbf05;
mem_array[23357] = 16'h6be4;
mem_array[23356] = 16'h3f5b;
mem_array[23359] = 16'h744d;
mem_array[23358] = 16'hbf1b;
mem_array[23361] = 16'habb8;
mem_array[23360] = 16'hbd7b;
mem_array[23363] = 16'h3474;
mem_array[23362] = 16'h3dec;
mem_array[23365] = 16'h6193;
mem_array[23364] = 16'h3dd1;
mem_array[23367] = 16'h3608;
mem_array[23366] = 16'h3f96;
mem_array[23369] = 16'h1836;
mem_array[23368] = 16'h3f11;
mem_array[23371] = 16'h7bc6;
mem_array[23370] = 16'h3f2d;
mem_array[23373] = 16'h16af;
mem_array[23372] = 16'hbf29;
mem_array[23375] = 16'h4604;
mem_array[23374] = 16'h3ec1;
mem_array[23377] = 16'h6028;
mem_array[23376] = 16'hbf57;
mem_array[23379] = 16'h2247;
mem_array[23378] = 16'h3ee1;
mem_array[23381] = 16'h2c56;
mem_array[23380] = 16'h3edd;
mem_array[23383] = 16'hbcef;
mem_array[23382] = 16'hbed8;
mem_array[23385] = 16'h2422;
mem_array[23384] = 16'hbf85;
mem_array[23387] = 16'hc356;
mem_array[23386] = 16'h3ea7;
mem_array[23389] = 16'h70e5;
mem_array[23388] = 16'h3ecc;
mem_array[23391] = 16'he6b2;
mem_array[23390] = 16'h3e6b;
mem_array[23393] = 16'hdfcd;
mem_array[23392] = 16'hbdb9;
mem_array[23395] = 16'h4f83;
mem_array[23394] = 16'h3c21;
mem_array[23397] = 16'h0997;
mem_array[23396] = 16'h3f82;
mem_array[23399] = 16'hcc3d;
mem_array[23398] = 16'hbe0b;
mem_array[23401] = 16'h71d4;
mem_array[23400] = 16'hbf7c;
mem_array[23403] = 16'hd168;
mem_array[23402] = 16'hbe98;
mem_array[23405] = 16'haab3;
mem_array[23404] = 16'h3f19;
mem_array[23407] = 16'h36a5;
mem_array[23406] = 16'hbf29;
mem_array[23409] = 16'h80de;
mem_array[23408] = 16'h3f18;
mem_array[23411] = 16'hf7b1;
mem_array[23410] = 16'hbe94;
mem_array[23413] = 16'hfcb1;
mem_array[23412] = 16'h3df5;
mem_array[23415] = 16'h094f;
mem_array[23414] = 16'h3e52;
mem_array[23417] = 16'hab49;
mem_array[23416] = 16'h3f2b;
mem_array[23419] = 16'h4749;
mem_array[23418] = 16'h3e36;
mem_array[23421] = 16'ha06f;
mem_array[23420] = 16'hbc90;
mem_array[23423] = 16'h1ff3;
mem_array[23422] = 16'h3dc7;
mem_array[23425] = 16'ha9e6;
mem_array[23424] = 16'hbe6e;
mem_array[23427] = 16'h8a26;
mem_array[23426] = 16'h3f0d;
mem_array[23429] = 16'h9bee;
mem_array[23428] = 16'h3dbf;
mem_array[23431] = 16'h7e99;
mem_array[23430] = 16'h3eea;
mem_array[23433] = 16'h9b7c;
mem_array[23432] = 16'h3e8d;
mem_array[23435] = 16'h8d9a;
mem_array[23434] = 16'hbae1;
mem_array[23437] = 16'h90b0;
mem_array[23436] = 16'hbee3;
mem_array[23439] = 16'hdae1;
mem_array[23438] = 16'h3dcf;
mem_array[23441] = 16'h6c2c;
mem_array[23440] = 16'h3edd;
mem_array[23443] = 16'h5326;
mem_array[23442] = 16'hbda1;
mem_array[23445] = 16'h36c3;
mem_array[23444] = 16'hbf91;
mem_array[23447] = 16'h1a8e;
mem_array[23446] = 16'hbdbc;
mem_array[23449] = 16'h3aaa;
mem_array[23448] = 16'h3f1a;
mem_array[23451] = 16'h623e;
mem_array[23450] = 16'hbe0a;
mem_array[23453] = 16'h2a4d;
mem_array[23452] = 16'h3e3d;
mem_array[23455] = 16'h525a;
mem_array[23454] = 16'hbd3e;
mem_array[23457] = 16'hc952;
mem_array[23456] = 16'h3fb1;
mem_array[23459] = 16'h0fe1;
mem_array[23458] = 16'h3d75;
mem_array[23461] = 16'h83b8;
mem_array[23460] = 16'h3d8a;
mem_array[23463] = 16'h85b4;
mem_array[23462] = 16'h3d0a;
mem_array[23465] = 16'h7304;
mem_array[23464] = 16'h3ee1;
mem_array[23467] = 16'ha303;
mem_array[23466] = 16'h3e29;
mem_array[23469] = 16'h4660;
mem_array[23468] = 16'h3d85;
mem_array[23471] = 16'h2592;
mem_array[23470] = 16'hbe0e;
mem_array[23473] = 16'hf216;
mem_array[23472] = 16'h3d1e;
mem_array[23475] = 16'he8dd;
mem_array[23474] = 16'h3ea2;
mem_array[23477] = 16'h2555;
mem_array[23476] = 16'h3ed3;
mem_array[23479] = 16'hb491;
mem_array[23478] = 16'h3d78;
mem_array[23481] = 16'h598e;
mem_array[23480] = 16'hbca2;
mem_array[23483] = 16'hbdf4;
mem_array[23482] = 16'hbda2;
mem_array[23485] = 16'h26ad;
mem_array[23484] = 16'h3e1b;
mem_array[23487] = 16'h9e6e;
mem_array[23486] = 16'h3e95;
mem_array[23489] = 16'hed49;
mem_array[23488] = 16'h3d5f;
mem_array[23491] = 16'hab7c;
mem_array[23490] = 16'hbe9c;
mem_array[23493] = 16'hf511;
mem_array[23492] = 16'h3e90;
mem_array[23495] = 16'h7337;
mem_array[23494] = 16'hbb72;
mem_array[23497] = 16'h895b;
mem_array[23496] = 16'hbe3c;
mem_array[23499] = 16'he51b;
mem_array[23498] = 16'hbd6c;
mem_array[23501] = 16'h1d91;
mem_array[23500] = 16'hbe48;
mem_array[23503] = 16'h9b84;
mem_array[23502] = 16'hbd05;
mem_array[23505] = 16'hf02e;
mem_array[23504] = 16'hbda9;
mem_array[23507] = 16'h8a1e;
mem_array[23506] = 16'h3d41;
mem_array[23509] = 16'h9270;
mem_array[23508] = 16'hbde8;
mem_array[23511] = 16'h3ef0;
mem_array[23510] = 16'h3d2c;
mem_array[23513] = 16'hcbdf;
mem_array[23512] = 16'h3df6;
mem_array[23515] = 16'h5d2d;
mem_array[23514] = 16'h3d2e;
mem_array[23517] = 16'h21cc;
mem_array[23516] = 16'h3f2d;
mem_array[23519] = 16'h05db;
mem_array[23518] = 16'hbe05;
mem_array[23521] = 16'h7d28;
mem_array[23520] = 16'h3da6;
mem_array[23523] = 16'h6d34;
mem_array[23522] = 16'hbc50;
mem_array[23525] = 16'h0f08;
mem_array[23524] = 16'h3cd9;
mem_array[23527] = 16'hdb6f;
mem_array[23526] = 16'hbd39;
mem_array[23529] = 16'h27db;
mem_array[23528] = 16'hbdca;
mem_array[23531] = 16'hcfd3;
mem_array[23530] = 16'h3f28;
mem_array[23533] = 16'h7f8e;
mem_array[23532] = 16'h3e84;
mem_array[23535] = 16'h338b;
mem_array[23534] = 16'hbcce;
mem_array[23537] = 16'h528c;
mem_array[23536] = 16'h3d8f;
mem_array[23539] = 16'h2534;
mem_array[23538] = 16'h3ad3;
mem_array[23541] = 16'h6fe4;
mem_array[23540] = 16'hbc23;
mem_array[23543] = 16'haf13;
mem_array[23542] = 16'h3d04;
mem_array[23545] = 16'ha0ac;
mem_array[23544] = 16'hbd8d;
mem_array[23547] = 16'he039;
mem_array[23546] = 16'hbd6f;
mem_array[23549] = 16'hd64b;
mem_array[23548] = 16'hbccd;
mem_array[23551] = 16'hc4e6;
mem_array[23550] = 16'hbea5;
mem_array[23553] = 16'h23a3;
mem_array[23552] = 16'h3d71;
mem_array[23555] = 16'h4094;
mem_array[23554] = 16'hbaa1;
mem_array[23557] = 16'ha705;
mem_array[23556] = 16'hbdb1;
mem_array[23559] = 16'hea8f;
mem_array[23558] = 16'hbda7;
mem_array[23561] = 16'h1720;
mem_array[23560] = 16'h3d86;
mem_array[23563] = 16'h9487;
mem_array[23562] = 16'h3f05;
mem_array[23565] = 16'hd899;
mem_array[23564] = 16'hbd73;
mem_array[23567] = 16'hf91d;
mem_array[23566] = 16'h3d40;
mem_array[23569] = 16'h8ca1;
mem_array[23568] = 16'hbd2c;
mem_array[23571] = 16'h986b;
mem_array[23570] = 16'hbdc9;
mem_array[23573] = 16'h3b68;
mem_array[23572] = 16'h3f74;
mem_array[23575] = 16'hce79;
mem_array[23574] = 16'hbcba;
mem_array[23577] = 16'h191e;
mem_array[23576] = 16'hbda6;
mem_array[23579] = 16'h58ec;
mem_array[23578] = 16'h3cbd;
mem_array[23581] = 16'hb0c4;
mem_array[23580] = 16'h3c9d;
mem_array[23583] = 16'h9f17;
mem_array[23582] = 16'h3e13;
mem_array[23585] = 16'h276e;
mem_array[23584] = 16'hbc2c;
mem_array[23587] = 16'h6f4b;
mem_array[23586] = 16'hbd87;
mem_array[23589] = 16'h682f;
mem_array[23588] = 16'h3d60;
mem_array[23591] = 16'he01d;
mem_array[23590] = 16'h3d13;
mem_array[23593] = 16'h40ef;
mem_array[23592] = 16'h3f0a;
mem_array[23595] = 16'h0c83;
mem_array[23594] = 16'h3e27;
mem_array[23597] = 16'h523e;
mem_array[23596] = 16'hbdac;
mem_array[23599] = 16'h4226;
mem_array[23598] = 16'hbbae;
mem_array[23601] = 16'h44c4;
mem_array[23600] = 16'h3cb7;
mem_array[23603] = 16'h411f;
mem_array[23602] = 16'h3db8;
mem_array[23605] = 16'h80dd;
mem_array[23604] = 16'hbe19;
mem_array[23607] = 16'he663;
mem_array[23606] = 16'hbeca;
mem_array[23609] = 16'hbf35;
mem_array[23608] = 16'hbd49;
mem_array[23611] = 16'hfd91;
mem_array[23610] = 16'hbebb;
mem_array[23613] = 16'h3b1f;
mem_array[23612] = 16'hbd9f;
mem_array[23615] = 16'hb6cf;
mem_array[23614] = 16'hbd28;
mem_array[23617] = 16'h34b3;
mem_array[23616] = 16'h3e96;
mem_array[23619] = 16'hc115;
mem_array[23618] = 16'h3e1f;
mem_array[23621] = 16'h30a6;
mem_array[23620] = 16'hbd08;
mem_array[23623] = 16'h90b8;
mem_array[23622] = 16'h3e05;
mem_array[23625] = 16'h13fc;
mem_array[23624] = 16'hbd03;
mem_array[23627] = 16'hd3f7;
mem_array[23626] = 16'hbe47;
mem_array[23629] = 16'hfa51;
mem_array[23628] = 16'h3f00;
mem_array[23631] = 16'h428e;
mem_array[23630] = 16'h3e1e;
mem_array[23633] = 16'h4ac3;
mem_array[23632] = 16'hbdec;
mem_array[23635] = 16'hd96c;
mem_array[23634] = 16'h3df7;
mem_array[23637] = 16'h9ddf;
mem_array[23636] = 16'hbd46;
mem_array[23639] = 16'hbf59;
mem_array[23638] = 16'hbc19;
mem_array[23641] = 16'hfca7;
mem_array[23640] = 16'h3ec2;
mem_array[23643] = 16'h66eb;
mem_array[23642] = 16'h3f95;
mem_array[23645] = 16'h194f;
mem_array[23644] = 16'h3d97;
mem_array[23647] = 16'h872e;
mem_array[23646] = 16'h3e0c;
mem_array[23649] = 16'hf72f;
mem_array[23648] = 16'hbd06;
mem_array[23651] = 16'hbaf0;
mem_array[23650] = 16'hbd74;
mem_array[23653] = 16'he120;
mem_array[23652] = 16'hbe83;
mem_array[23655] = 16'h08ff;
mem_array[23654] = 16'h3f2c;
mem_array[23657] = 16'h08b5;
mem_array[23656] = 16'hbe46;
mem_array[23659] = 16'h8af3;
mem_array[23658] = 16'hbd2f;
mem_array[23661] = 16'hdf92;
mem_array[23660] = 16'h3ca5;
mem_array[23663] = 16'hf6ff;
mem_array[23662] = 16'hbdd3;
mem_array[23665] = 16'ha34a;
mem_array[23664] = 16'h3ec6;
mem_array[23667] = 16'ha595;
mem_array[23666] = 16'hbf59;
mem_array[23669] = 16'hff92;
mem_array[23668] = 16'hbdd6;
mem_array[23671] = 16'hd04c;
mem_array[23670] = 16'hbeee;
mem_array[23673] = 16'h93f2;
mem_array[23672] = 16'h3f1d;
mem_array[23675] = 16'h4548;
mem_array[23674] = 16'hbed0;
mem_array[23677] = 16'hf1f0;
mem_array[23676] = 16'hbe4e;
mem_array[23679] = 16'h2613;
mem_array[23678] = 16'hbe0e;
mem_array[23681] = 16'hdd32;
mem_array[23680] = 16'hbe64;
mem_array[23683] = 16'h9613;
mem_array[23682] = 16'h3f46;
mem_array[23685] = 16'h09ad;
mem_array[23684] = 16'h3d86;
mem_array[23687] = 16'h8fe6;
mem_array[23686] = 16'hbeb4;
mem_array[23689] = 16'hffdc;
mem_array[23688] = 16'hbf10;
mem_array[23691] = 16'hcedf;
mem_array[23690] = 16'h3f21;
mem_array[23693] = 16'h8caf;
mem_array[23692] = 16'h3ef0;
mem_array[23695] = 16'h0532;
mem_array[23694] = 16'h3f2e;
mem_array[23697] = 16'h9210;
mem_array[23696] = 16'hbf05;
mem_array[23699] = 16'hc3d2;
mem_array[23698] = 16'hbf2f;
mem_array[23701] = 16'h3f54;
mem_array[23700] = 16'h3ea0;
mem_array[23703] = 16'h2028;
mem_array[23702] = 16'h3ebc;
mem_array[23705] = 16'h4318;
mem_array[23704] = 16'h3f0a;
mem_array[23707] = 16'h3ae9;
mem_array[23706] = 16'hbf25;
mem_array[23709] = 16'hb5eb;
mem_array[23708] = 16'hbd9a;
mem_array[23711] = 16'he89d;
mem_array[23710] = 16'h3d1a;
mem_array[23713] = 16'h2c5c;
mem_array[23712] = 16'h3e43;
mem_array[23715] = 16'he370;
mem_array[23714] = 16'h3f43;
mem_array[23717] = 16'he2ca;
mem_array[23716] = 16'hbf67;
mem_array[23719] = 16'h3dda;
mem_array[23718] = 16'hbe41;
mem_array[23721] = 16'h1e9b;
mem_array[23720] = 16'h3ccf;
mem_array[23723] = 16'h7ebf;
mem_array[23722] = 16'h3d3b;
mem_array[23725] = 16'hfe7a;
mem_array[23724] = 16'hbf82;
mem_array[23727] = 16'hddba;
mem_array[23726] = 16'hbdd2;
mem_array[23729] = 16'hfbf3;
mem_array[23728] = 16'hbf1f;
mem_array[23731] = 16'h01b6;
mem_array[23730] = 16'h3f1e;
mem_array[23733] = 16'hf543;
mem_array[23732] = 16'h3f08;
mem_array[23735] = 16'h9166;
mem_array[23734] = 16'h3e7d;
mem_array[23737] = 16'h5425;
mem_array[23736] = 16'h3e1e;
mem_array[23739] = 16'h1635;
mem_array[23738] = 16'hbf1c;
mem_array[23741] = 16'hbd18;
mem_array[23740] = 16'hbf8a;
mem_array[23743] = 16'h2e3a;
mem_array[23742] = 16'hbf08;
mem_array[23745] = 16'h2c68;
mem_array[23744] = 16'hbe92;
mem_array[23747] = 16'h6a51;
mem_array[23746] = 16'hbe5c;
mem_array[23749] = 16'hdac5;
mem_array[23748] = 16'hbf93;
mem_array[23751] = 16'h9489;
mem_array[23750] = 16'h3f11;
mem_array[23753] = 16'hf101;
mem_array[23752] = 16'h3dfb;
mem_array[23755] = 16'h2bf3;
mem_array[23754] = 16'hbcae;
mem_array[23757] = 16'h9465;
mem_array[23756] = 16'h3f0f;
mem_array[23759] = 16'h66e2;
mem_array[23758] = 16'h3dc7;
mem_array[23761] = 16'hf4ed;
mem_array[23760] = 16'hbdf0;
mem_array[23763] = 16'h2abc;
mem_array[23762] = 16'hbebd;
mem_array[23765] = 16'h9f28;
mem_array[23764] = 16'hbeec;
mem_array[23767] = 16'he727;
mem_array[23766] = 16'hbee1;
mem_array[23769] = 16'hd790;
mem_array[23768] = 16'h3d26;
mem_array[23771] = 16'hb166;
mem_array[23770] = 16'hbe59;
mem_array[23773] = 16'h98f0;
mem_array[23772] = 16'hbd2c;
mem_array[23775] = 16'h44fc;
mem_array[23774] = 16'h3f27;
mem_array[23777] = 16'h1cd0;
mem_array[23776] = 16'hbf93;
mem_array[23779] = 16'habe1;
mem_array[23778] = 16'h3f65;
mem_array[23781] = 16'h78e9;
mem_array[23780] = 16'hbd98;
mem_array[23783] = 16'ha803;
mem_array[23782] = 16'hbd48;
mem_array[23785] = 16'h393f;
mem_array[23784] = 16'hbe25;
mem_array[23787] = 16'ha071;
mem_array[23786] = 16'h3e74;
mem_array[23789] = 16'had0a;
mem_array[23788] = 16'hbea8;
mem_array[23791] = 16'h52d7;
mem_array[23790] = 16'h3ef1;
mem_array[23793] = 16'h1748;
mem_array[23792] = 16'hbe89;
mem_array[23795] = 16'h4a72;
mem_array[23794] = 16'hbe29;
mem_array[23797] = 16'h85da;
mem_array[23796] = 16'h3eef;
mem_array[23799] = 16'he6f5;
mem_array[23798] = 16'hbe85;
mem_array[23801] = 16'hef58;
mem_array[23800] = 16'hbf42;
mem_array[23803] = 16'h92ae;
mem_array[23802] = 16'h3ea4;
mem_array[23805] = 16'hd913;
mem_array[23804] = 16'hbe61;
mem_array[23807] = 16'hac46;
mem_array[23806] = 16'h3ea1;
mem_array[23809] = 16'h77bc;
mem_array[23808] = 16'hbfcd;
mem_array[23811] = 16'heb35;
mem_array[23810] = 16'hbe9f;
mem_array[23813] = 16'hb45a;
mem_array[23812] = 16'hbe54;
mem_array[23815] = 16'h3cc3;
mem_array[23814] = 16'hbd46;
mem_array[23817] = 16'hcdfb;
mem_array[23816] = 16'hbe32;
mem_array[23819] = 16'h5a2d;
mem_array[23818] = 16'h3f06;
mem_array[23821] = 16'h3095;
mem_array[23820] = 16'hbf16;
mem_array[23823] = 16'h201d;
mem_array[23822] = 16'hbce8;
mem_array[23825] = 16'hc78e;
mem_array[23824] = 16'hbf23;
mem_array[23827] = 16'h14c4;
mem_array[23826] = 16'h3e4f;
mem_array[23829] = 16'hb63d;
mem_array[23828] = 16'h3c36;
mem_array[23831] = 16'hff6c;
mem_array[23830] = 16'hbeab;
mem_array[23833] = 16'hdf77;
mem_array[23832] = 16'hbe94;
mem_array[23835] = 16'h60da;
mem_array[23834] = 16'h3ee2;
mem_array[23837] = 16'hdcad;
mem_array[23836] = 16'hbf81;
mem_array[23839] = 16'h4efa;
mem_array[23838] = 16'h3dd6;
mem_array[23841] = 16'h6b45;
mem_array[23840] = 16'hbc8f;
mem_array[23843] = 16'h3aca;
mem_array[23842] = 16'h3d2e;
mem_array[23845] = 16'hbe7d;
mem_array[23844] = 16'h3e6b;
mem_array[23847] = 16'hea12;
mem_array[23846] = 16'hbf3d;
mem_array[23849] = 16'h61b4;
mem_array[23848] = 16'hbf7f;
mem_array[23851] = 16'hc02d;
mem_array[23850] = 16'hbe86;
mem_array[23853] = 16'h3f0a;
mem_array[23852] = 16'hbfa1;
mem_array[23855] = 16'ha6fa;
mem_array[23854] = 16'h3f35;
mem_array[23857] = 16'hf87f;
mem_array[23856] = 16'h3e34;
mem_array[23859] = 16'hc792;
mem_array[23858] = 16'h3e51;
mem_array[23861] = 16'he8a2;
mem_array[23860] = 16'hbd22;
mem_array[23863] = 16'h0b9b;
mem_array[23862] = 16'h3daa;
mem_array[23865] = 16'h5d4f;
mem_array[23864] = 16'h3e83;
mem_array[23867] = 16'h0e5b;
mem_array[23866] = 16'h3ce8;
mem_array[23869] = 16'h14de;
mem_array[23868] = 16'hbf80;
mem_array[23871] = 16'h7680;
mem_array[23870] = 16'h3ef0;
mem_array[23873] = 16'h6a45;
mem_array[23872] = 16'hbeef;
mem_array[23875] = 16'h432d;
mem_array[23874] = 16'h3edb;
mem_array[23877] = 16'hfef9;
mem_array[23876] = 16'h3edf;
mem_array[23879] = 16'h464b;
mem_array[23878] = 16'h3f0a;
mem_array[23881] = 16'h9cd9;
mem_array[23880] = 16'hbec1;
mem_array[23883] = 16'he914;
mem_array[23882] = 16'hbd26;
mem_array[23885] = 16'h6251;
mem_array[23884] = 16'h3f03;
mem_array[23887] = 16'hd583;
mem_array[23886] = 16'h3f07;
mem_array[23889] = 16'hb253;
mem_array[23888] = 16'h3df3;
mem_array[23891] = 16'h1bdf;
mem_array[23890] = 16'hbe96;
mem_array[23893] = 16'haff7;
mem_array[23892] = 16'h3e64;
mem_array[23895] = 16'hf0ef;
mem_array[23894] = 16'hbebd;
mem_array[23897] = 16'hc2b5;
mem_array[23896] = 16'hc001;
mem_array[23899] = 16'hed27;
mem_array[23898] = 16'hbe8f;
mem_array[23901] = 16'h07b5;
mem_array[23900] = 16'hbb96;
mem_array[23903] = 16'h2a56;
mem_array[23902] = 16'hbdc9;
mem_array[23905] = 16'h84aa;
mem_array[23904] = 16'h3e5d;
mem_array[23907] = 16'h2693;
mem_array[23906] = 16'h3e93;
mem_array[23909] = 16'h2b2b;
mem_array[23908] = 16'hbfa1;
mem_array[23911] = 16'h4238;
mem_array[23910] = 16'hbeb3;
mem_array[23913] = 16'h9576;
mem_array[23912] = 16'hbfcb;
mem_array[23915] = 16'h9c6d;
mem_array[23914] = 16'h3db5;
mem_array[23917] = 16'hbdf3;
mem_array[23916] = 16'hbe70;
mem_array[23919] = 16'h0fa8;
mem_array[23918] = 16'hbe24;
mem_array[23921] = 16'h7259;
mem_array[23920] = 16'hbbf0;
mem_array[23923] = 16'h88f6;
mem_array[23922] = 16'h3eb7;
mem_array[23925] = 16'h331f;
mem_array[23924] = 16'h3e4f;
mem_array[23927] = 16'hd4cc;
mem_array[23926] = 16'h3e97;
mem_array[23929] = 16'h54bf;
mem_array[23928] = 16'hbfa6;
mem_array[23931] = 16'h4cb4;
mem_array[23930] = 16'h3ccc;
mem_array[23933] = 16'h5b7b;
mem_array[23932] = 16'hbe44;
mem_array[23935] = 16'hb77c;
mem_array[23934] = 16'h3e0f;
mem_array[23937] = 16'h1e67;
mem_array[23936] = 16'h3f50;
mem_array[23939] = 16'h6a43;
mem_array[23938] = 16'h3eb2;
mem_array[23941] = 16'h2ac8;
mem_array[23940] = 16'h3eec;
mem_array[23943] = 16'had6c;
mem_array[23942] = 16'hbe9c;
mem_array[23945] = 16'hecd6;
mem_array[23944] = 16'hbdc2;
mem_array[23947] = 16'h4f10;
mem_array[23946] = 16'h3edc;
mem_array[23949] = 16'h82d8;
mem_array[23948] = 16'h3e95;
mem_array[23951] = 16'h4afc;
mem_array[23950] = 16'hbe3d;
mem_array[23953] = 16'he484;
mem_array[23952] = 16'h3df0;
mem_array[23955] = 16'h7bff;
mem_array[23954] = 16'hbf04;
mem_array[23957] = 16'h3cbe;
mem_array[23956] = 16'hbf99;
mem_array[23959] = 16'h61ea;
mem_array[23958] = 16'hbd28;
mem_array[23961] = 16'hf3c3;
mem_array[23960] = 16'hbc5c;
mem_array[23963] = 16'hb4ab;
mem_array[23962] = 16'hbac2;
mem_array[23965] = 16'h0396;
mem_array[23964] = 16'h3e02;
mem_array[23967] = 16'ha281;
mem_array[23966] = 16'h3efc;
mem_array[23969] = 16'h8f93;
mem_array[23968] = 16'hbf8f;
mem_array[23971] = 16'hfff8;
mem_array[23970] = 16'hbe21;
mem_array[23973] = 16'h63e2;
mem_array[23972] = 16'hbf67;
mem_array[23975] = 16'he173;
mem_array[23974] = 16'h3ec0;
mem_array[23977] = 16'ha415;
mem_array[23976] = 16'h3d67;
mem_array[23979] = 16'h9e57;
mem_array[23978] = 16'h3d97;
mem_array[23981] = 16'he9e3;
mem_array[23980] = 16'h3e90;
mem_array[23983] = 16'h55e4;
mem_array[23982] = 16'h3de6;
mem_array[23985] = 16'h4c94;
mem_array[23984] = 16'h3f01;
mem_array[23987] = 16'h4d27;
mem_array[23986] = 16'h3e95;
mem_array[23989] = 16'he3f5;
mem_array[23988] = 16'hbe3c;
mem_array[23991] = 16'h6330;
mem_array[23990] = 16'h3e3c;
mem_array[23993] = 16'h4709;
mem_array[23992] = 16'hbdf5;
mem_array[23995] = 16'h6aaf;
mem_array[23994] = 16'hbc74;
mem_array[23997] = 16'h582f;
mem_array[23996] = 16'h3f3f;
mem_array[23999] = 16'h816f;
mem_array[23998] = 16'h3e5d;
mem_array[24001] = 16'h3611;
mem_array[24000] = 16'h3e5e;
mem_array[24003] = 16'hc60a;
mem_array[24002] = 16'hbbf0;
mem_array[24005] = 16'h68fa;
mem_array[24004] = 16'hbfc0;
mem_array[24007] = 16'ha888;
mem_array[24006] = 16'h3ecd;
mem_array[24009] = 16'h5eec;
mem_array[24008] = 16'hbdab;
mem_array[24011] = 16'hcffb;
mem_array[24010] = 16'hbe20;
mem_array[24013] = 16'h321e;
mem_array[24012] = 16'hbc50;
mem_array[24015] = 16'he900;
mem_array[24014] = 16'hbdc8;
mem_array[24017] = 16'h1fd8;
mem_array[24016] = 16'hbf8f;
mem_array[24019] = 16'h86b1;
mem_array[24018] = 16'h3f4a;
mem_array[24021] = 16'hacf6;
mem_array[24020] = 16'hbc42;
mem_array[24023] = 16'hafca;
mem_array[24022] = 16'h3c82;
mem_array[24025] = 16'had60;
mem_array[24024] = 16'h3e9f;
mem_array[24027] = 16'h6a9c;
mem_array[24026] = 16'h3ebc;
mem_array[24029] = 16'h5a45;
mem_array[24028] = 16'hbfd1;
mem_array[24031] = 16'h90c3;
mem_array[24030] = 16'hbdcb;
mem_array[24033] = 16'h01cf;
mem_array[24032] = 16'hbebb;
mem_array[24035] = 16'h2595;
mem_array[24034] = 16'h3e16;
mem_array[24037] = 16'h7198;
mem_array[24036] = 16'hbe11;
mem_array[24039] = 16'h00fa;
mem_array[24038] = 16'h3d29;
mem_array[24041] = 16'h0200;
mem_array[24040] = 16'h3e53;
mem_array[24043] = 16'h08fa;
mem_array[24042] = 16'h3e53;
mem_array[24045] = 16'h1c8d;
mem_array[24044] = 16'h3f22;
mem_array[24047] = 16'he9de;
mem_array[24046] = 16'h3e5c;
mem_array[24049] = 16'h1725;
mem_array[24048] = 16'h3e48;
mem_array[24051] = 16'h165b;
mem_array[24050] = 16'h3b49;
mem_array[24053] = 16'h5b35;
mem_array[24052] = 16'hbd87;
mem_array[24055] = 16'h4903;
mem_array[24054] = 16'h3d34;
mem_array[24057] = 16'h8d5b;
mem_array[24056] = 16'h3e83;
mem_array[24059] = 16'hc883;
mem_array[24058] = 16'h3e94;
mem_array[24061] = 16'h074f;
mem_array[24060] = 16'hbed2;
mem_array[24063] = 16'h82ce;
mem_array[24062] = 16'h3e22;
mem_array[24065] = 16'ha503;
mem_array[24064] = 16'hc002;
mem_array[24067] = 16'h1678;
mem_array[24066] = 16'h3e1b;
mem_array[24069] = 16'h1491;
mem_array[24068] = 16'h3e18;
mem_array[24071] = 16'h2588;
mem_array[24070] = 16'hbdd7;
mem_array[24073] = 16'h0599;
mem_array[24072] = 16'hbe9b;
mem_array[24075] = 16'ha816;
mem_array[24074] = 16'hbc18;
mem_array[24077] = 16'h6f45;
mem_array[24076] = 16'hbf4f;
mem_array[24079] = 16'h2cdc;
mem_array[24078] = 16'h3de0;
mem_array[24081] = 16'h0dea;
mem_array[24080] = 16'hbcd5;
mem_array[24083] = 16'h6b93;
mem_array[24082] = 16'hbd5d;
mem_array[24085] = 16'h301d;
mem_array[24084] = 16'h3dda;
mem_array[24087] = 16'h7f77;
mem_array[24086] = 16'h3f40;
mem_array[24089] = 16'h2686;
mem_array[24088] = 16'hbfb9;
mem_array[24091] = 16'h7194;
mem_array[24090] = 16'hbd30;
mem_array[24093] = 16'h6f79;
mem_array[24092] = 16'hbf56;
mem_array[24095] = 16'hbe18;
mem_array[24094] = 16'h3ec5;
mem_array[24097] = 16'h95b5;
mem_array[24096] = 16'hbd70;
mem_array[24099] = 16'h7b66;
mem_array[24098] = 16'h3e86;
mem_array[24101] = 16'he2b2;
mem_array[24100] = 16'h3e54;
mem_array[24103] = 16'h8407;
mem_array[24102] = 16'h3e93;
mem_array[24105] = 16'h74a5;
mem_array[24104] = 16'h3dcc;
mem_array[24107] = 16'hcde8;
mem_array[24106] = 16'h3de1;
mem_array[24109] = 16'h07e4;
mem_array[24108] = 16'h3e3c;
mem_array[24111] = 16'hf497;
mem_array[24110] = 16'h3d33;
mem_array[24113] = 16'h8018;
mem_array[24112] = 16'hbea1;
mem_array[24115] = 16'h30eb;
mem_array[24114] = 16'h3dec;
mem_array[24117] = 16'h0b28;
mem_array[24116] = 16'h3e78;
mem_array[24119] = 16'h28f1;
mem_array[24118] = 16'h3ed2;
mem_array[24121] = 16'h9fd2;
mem_array[24120] = 16'hbec2;
mem_array[24123] = 16'hbbc1;
mem_array[24122] = 16'h3dd5;
mem_array[24125] = 16'h8344;
mem_array[24124] = 16'hc006;
mem_array[24127] = 16'hd593;
mem_array[24126] = 16'h3e26;
mem_array[24129] = 16'h1eed;
mem_array[24128] = 16'hbea9;
mem_array[24131] = 16'h7109;
mem_array[24130] = 16'h3e5c;
mem_array[24133] = 16'ha0bf;
mem_array[24132] = 16'hbe84;
mem_array[24135] = 16'hb7b0;
mem_array[24134] = 16'hbd88;
mem_array[24137] = 16'hf2b6;
mem_array[24136] = 16'hbd38;
mem_array[24139] = 16'h16d9;
mem_array[24138] = 16'hbf67;
mem_array[24141] = 16'hd2da;
mem_array[24140] = 16'hbd95;
mem_array[24143] = 16'h95b4;
mem_array[24142] = 16'hbdb5;
mem_array[24145] = 16'hb3e4;
mem_array[24144] = 16'hbd2d;
mem_array[24147] = 16'h8cd5;
mem_array[24146] = 16'h3dc1;
mem_array[24149] = 16'hc46d;
mem_array[24148] = 16'hbfc0;
mem_array[24151] = 16'hc4a1;
mem_array[24150] = 16'hbae7;
mem_array[24153] = 16'hc786;
mem_array[24152] = 16'hbe7d;
mem_array[24155] = 16'h17f2;
mem_array[24154] = 16'h3e92;
mem_array[24157] = 16'ha205;
mem_array[24156] = 16'h3dd3;
mem_array[24159] = 16'hf1d5;
mem_array[24158] = 16'h3d30;
mem_array[24161] = 16'h74de;
mem_array[24160] = 16'hbd25;
mem_array[24163] = 16'h6c52;
mem_array[24162] = 16'h3e13;
mem_array[24165] = 16'he055;
mem_array[24164] = 16'h3e16;
mem_array[24167] = 16'ha013;
mem_array[24166] = 16'h3dd8;
mem_array[24169] = 16'h8b63;
mem_array[24168] = 16'h3dca;
mem_array[24171] = 16'h0d12;
mem_array[24170] = 16'hbe9d;
mem_array[24173] = 16'h61fe;
mem_array[24172] = 16'hbd72;
mem_array[24175] = 16'h495e;
mem_array[24174] = 16'h3e1f;
mem_array[24177] = 16'hb2cb;
mem_array[24176] = 16'h3ec6;
mem_array[24179] = 16'h0cb6;
mem_array[24178] = 16'h3ed3;
mem_array[24181] = 16'h43ec;
mem_array[24180] = 16'h3ce2;
mem_array[24183] = 16'h1e3e;
mem_array[24182] = 16'h3e9a;
mem_array[24185] = 16'h129d;
mem_array[24184] = 16'hbefa;
mem_array[24187] = 16'h2988;
mem_array[24186] = 16'h3dec;
mem_array[24189] = 16'h14cf;
mem_array[24188] = 16'hbe47;
mem_array[24191] = 16'he607;
mem_array[24190] = 16'hbdeb;
mem_array[24193] = 16'hd9f2;
mem_array[24192] = 16'hbe7a;
mem_array[24195] = 16'h39c2;
mem_array[24194] = 16'hbbe4;
mem_array[24197] = 16'h13f0;
mem_array[24196] = 16'hbd02;
mem_array[24199] = 16'h1b8d;
mem_array[24198] = 16'hbeb5;
mem_array[24201] = 16'h8b83;
mem_array[24200] = 16'hbca4;
mem_array[24203] = 16'hd4c2;
mem_array[24202] = 16'h3cc2;
mem_array[24205] = 16'h5519;
mem_array[24204] = 16'h3d46;
mem_array[24207] = 16'hfb16;
mem_array[24206] = 16'h3e79;
mem_array[24209] = 16'hc869;
mem_array[24208] = 16'hbed4;
mem_array[24211] = 16'h3201;
mem_array[24210] = 16'h3daa;
mem_array[24213] = 16'h295c;
mem_array[24212] = 16'hbe0f;
mem_array[24215] = 16'h6d5e;
mem_array[24214] = 16'h3e46;
mem_array[24217] = 16'h58ba;
mem_array[24216] = 16'h3d87;
mem_array[24219] = 16'h4548;
mem_array[24218] = 16'h3db3;
mem_array[24221] = 16'h6e0b;
mem_array[24220] = 16'h3ea1;
mem_array[24223] = 16'h3850;
mem_array[24222] = 16'hbbe4;
mem_array[24225] = 16'hd310;
mem_array[24224] = 16'hbdc6;
mem_array[24227] = 16'hd64a;
mem_array[24226] = 16'h3e13;
mem_array[24229] = 16'h98a5;
mem_array[24228] = 16'h3ea0;
mem_array[24231] = 16'h6993;
mem_array[24230] = 16'hbf20;
mem_array[24233] = 16'he45b;
mem_array[24232] = 16'h3e11;
mem_array[24235] = 16'h3585;
mem_array[24234] = 16'h3e19;
mem_array[24237] = 16'hd4da;
mem_array[24236] = 16'h3ee0;
mem_array[24239] = 16'h9b64;
mem_array[24238] = 16'h3f24;
mem_array[24241] = 16'h8c3f;
mem_array[24240] = 16'hbe3c;
mem_array[24243] = 16'h52ab;
mem_array[24242] = 16'hbe74;
mem_array[24245] = 16'h31de;
mem_array[24244] = 16'hbe12;
mem_array[24247] = 16'hefc3;
mem_array[24246] = 16'hbecf;
mem_array[24249] = 16'h6549;
mem_array[24248] = 16'hbea8;
mem_array[24251] = 16'h3e7d;
mem_array[24250] = 16'h3d8b;
mem_array[24253] = 16'h5e67;
mem_array[24252] = 16'hbd92;
mem_array[24255] = 16'h844b;
mem_array[24254] = 16'h3db0;
mem_array[24257] = 16'ha37e;
mem_array[24256] = 16'hbdce;
mem_array[24259] = 16'hc312;
mem_array[24258] = 16'hbe85;
mem_array[24261] = 16'h38f4;
mem_array[24260] = 16'h3d9d;
mem_array[24263] = 16'hac71;
mem_array[24262] = 16'hbd8f;
mem_array[24265] = 16'he4d6;
mem_array[24264] = 16'h3e43;
mem_array[24267] = 16'h1ac4;
mem_array[24266] = 16'h3ed5;
mem_array[24269] = 16'h4bb8;
mem_array[24268] = 16'hbe86;
mem_array[24271] = 16'hb269;
mem_array[24270] = 16'h3e2f;
mem_array[24273] = 16'h2038;
mem_array[24272] = 16'hbe76;
mem_array[24275] = 16'h4e64;
mem_array[24274] = 16'hbe0b;
mem_array[24277] = 16'hdd48;
mem_array[24276] = 16'hbe46;
mem_array[24279] = 16'hcca5;
mem_array[24278] = 16'hbd8f;
mem_array[24281] = 16'hdf39;
mem_array[24280] = 16'h3e5d;
mem_array[24283] = 16'haa37;
mem_array[24282] = 16'hbcbb;
mem_array[24285] = 16'ha09e;
mem_array[24284] = 16'h3ec9;
mem_array[24287] = 16'h493c;
mem_array[24286] = 16'h3e48;
mem_array[24289] = 16'h616e;
mem_array[24288] = 16'h3e4f;
mem_array[24291] = 16'h3b5c;
mem_array[24290] = 16'hbf4c;
mem_array[24293] = 16'h4fb9;
mem_array[24292] = 16'h3de7;
mem_array[24295] = 16'ha132;
mem_array[24294] = 16'h3cae;
mem_array[24297] = 16'h912c;
mem_array[24296] = 16'h3e2d;
mem_array[24299] = 16'haf78;
mem_array[24298] = 16'h3dae;
mem_array[24301] = 16'hd472;
mem_array[24300] = 16'h3e08;
mem_array[24303] = 16'he786;
mem_array[24302] = 16'hc001;
mem_array[24305] = 16'h73c1;
mem_array[24304] = 16'hbe1c;
mem_array[24307] = 16'h1fb2;
mem_array[24306] = 16'hbf48;
mem_array[24309] = 16'hab15;
mem_array[24308] = 16'hbde9;
mem_array[24311] = 16'h37da;
mem_array[24310] = 16'h3d94;
mem_array[24313] = 16'hde12;
mem_array[24312] = 16'hbd93;
mem_array[24315] = 16'ha152;
mem_array[24314] = 16'h3d9f;
mem_array[24317] = 16'he46b;
mem_array[24316] = 16'hbd87;
mem_array[24319] = 16'h09ff;
mem_array[24318] = 16'hbe92;
mem_array[24321] = 16'h2cd0;
mem_array[24320] = 16'hbd0b;
mem_array[24323] = 16'h4e20;
mem_array[24322] = 16'hbb97;
mem_array[24325] = 16'h28d4;
mem_array[24324] = 16'h3e2a;
mem_array[24327] = 16'h6ac1;
mem_array[24326] = 16'h3e41;
mem_array[24329] = 16'h5fdb;
mem_array[24328] = 16'hbf5f;
mem_array[24331] = 16'h5eff;
mem_array[24330] = 16'h3e85;
mem_array[24333] = 16'h4092;
mem_array[24332] = 16'h3d15;
mem_array[24335] = 16'h4870;
mem_array[24334] = 16'hbe2a;
mem_array[24337] = 16'h4572;
mem_array[24336] = 16'h3d9b;
mem_array[24339] = 16'h0ab6;
mem_array[24338] = 16'hbebf;
mem_array[24341] = 16'h81b9;
mem_array[24340] = 16'h3d73;
mem_array[24343] = 16'haf82;
mem_array[24342] = 16'h3d5c;
mem_array[24345] = 16'h6e0d;
mem_array[24344] = 16'hbdc5;
mem_array[24347] = 16'h77b8;
mem_array[24346] = 16'h3d27;
mem_array[24349] = 16'h2320;
mem_array[24348] = 16'h3e3a;
mem_array[24351] = 16'h3488;
mem_array[24350] = 16'hbfc5;
mem_array[24353] = 16'h95f3;
mem_array[24352] = 16'hbd92;
mem_array[24355] = 16'h9b2a;
mem_array[24354] = 16'hbd2d;
mem_array[24357] = 16'h3c5f;
mem_array[24356] = 16'h3de8;
mem_array[24359] = 16'h4cf0;
mem_array[24358] = 16'hbe9d;
mem_array[24361] = 16'h6eba;
mem_array[24360] = 16'h3e68;
mem_array[24363] = 16'hded4;
mem_array[24362] = 16'hbf80;
mem_array[24365] = 16'h2641;
mem_array[24364] = 16'hbe3e;
mem_array[24367] = 16'he237;
mem_array[24366] = 16'hbf86;
mem_array[24369] = 16'h2f4c;
mem_array[24368] = 16'h3e43;
mem_array[24371] = 16'ha373;
mem_array[24370] = 16'h3e3b;
mem_array[24373] = 16'h469d;
mem_array[24372] = 16'h3eb2;
mem_array[24375] = 16'h5198;
mem_array[24374] = 16'h3cab;
mem_array[24377] = 16'hf90c;
mem_array[24376] = 16'hbe55;
mem_array[24379] = 16'h3192;
mem_array[24378] = 16'h3ea2;
mem_array[24381] = 16'heff9;
mem_array[24380] = 16'hbd59;
mem_array[24383] = 16'h09fc;
mem_array[24382] = 16'hbcd1;
mem_array[24385] = 16'hd420;
mem_array[24384] = 16'hbd6b;
mem_array[24387] = 16'h86cd;
mem_array[24386] = 16'h3e39;
mem_array[24389] = 16'h8469;
mem_array[24388] = 16'hbf55;
mem_array[24391] = 16'h1017;
mem_array[24390] = 16'h3e87;
mem_array[24393] = 16'h8c0f;
mem_array[24392] = 16'h3dc9;
mem_array[24395] = 16'he1eb;
mem_array[24394] = 16'h3dbb;
mem_array[24397] = 16'h762d;
mem_array[24396] = 16'h3dd0;
mem_array[24399] = 16'h3860;
mem_array[24398] = 16'hbf08;
mem_array[24401] = 16'he650;
mem_array[24400] = 16'hbd4c;
mem_array[24403] = 16'h22a4;
mem_array[24402] = 16'h3cfe;
mem_array[24405] = 16'h9e78;
mem_array[24404] = 16'hbea6;
mem_array[24407] = 16'hb458;
mem_array[24406] = 16'hbe07;
mem_array[24409] = 16'ha802;
mem_array[24408] = 16'h3eea;
mem_array[24411] = 16'had66;
mem_array[24410] = 16'hbe75;
mem_array[24413] = 16'hfb35;
mem_array[24412] = 16'hbd73;
mem_array[24415] = 16'he354;
mem_array[24414] = 16'hbe8c;
mem_array[24417] = 16'h7a8a;
mem_array[24416] = 16'hbd4d;
mem_array[24419] = 16'h3566;
mem_array[24418] = 16'hbf17;
mem_array[24421] = 16'haae7;
mem_array[24420] = 16'hbd67;
mem_array[24423] = 16'he64d;
mem_array[24422] = 16'hbed8;
mem_array[24425] = 16'ha86c;
mem_array[24424] = 16'hbe73;
mem_array[24427] = 16'h0aaa;
mem_array[24426] = 16'hbf81;
mem_array[24429] = 16'h3302;
mem_array[24428] = 16'h3eb3;
mem_array[24431] = 16'h4ce9;
mem_array[24430] = 16'h3d24;
mem_array[24433] = 16'h2900;
mem_array[24432] = 16'h3e8b;
mem_array[24435] = 16'h78d2;
mem_array[24434] = 16'hbc05;
mem_array[24437] = 16'hc5e9;
mem_array[24436] = 16'hbe42;
mem_array[24439] = 16'hd881;
mem_array[24438] = 16'hbd18;
mem_array[24441] = 16'hc435;
mem_array[24440] = 16'hbcb7;
mem_array[24443] = 16'h30b8;
mem_array[24442] = 16'hbd9e;
mem_array[24445] = 16'h03e1;
mem_array[24444] = 16'hbd91;
mem_array[24447] = 16'h1fe5;
mem_array[24446] = 16'hbe8b;
mem_array[24449] = 16'h53dd;
mem_array[24448] = 16'hbdfe;
mem_array[24451] = 16'h3608;
mem_array[24450] = 16'h3e72;
mem_array[24453] = 16'h1372;
mem_array[24452] = 16'hbc55;
mem_array[24455] = 16'h11a7;
mem_array[24454] = 16'hbd85;
mem_array[24457] = 16'hf680;
mem_array[24456] = 16'h3e05;
mem_array[24459] = 16'hf175;
mem_array[24458] = 16'hbf27;
mem_array[24461] = 16'h20cf;
mem_array[24460] = 16'h3e6d;
mem_array[24463] = 16'h7d28;
mem_array[24462] = 16'h3dfe;
mem_array[24465] = 16'h6b34;
mem_array[24464] = 16'hbe92;
mem_array[24467] = 16'hc115;
mem_array[24466] = 16'hbe46;
mem_array[24469] = 16'h7104;
mem_array[24468] = 16'h3d5a;
mem_array[24471] = 16'h135a;
mem_array[24470] = 16'h3d8c;
mem_array[24473] = 16'hc234;
mem_array[24472] = 16'hbb8b;
mem_array[24475] = 16'hb9df;
mem_array[24474] = 16'hbd94;
mem_array[24477] = 16'he28f;
mem_array[24476] = 16'h3e2a;
mem_array[24479] = 16'hbb38;
mem_array[24478] = 16'hbe94;
mem_array[24481] = 16'he02d;
mem_array[24480] = 16'h3ddc;
mem_array[24483] = 16'h2ece;
mem_array[24482] = 16'h3d76;
mem_array[24485] = 16'hb244;
mem_array[24484] = 16'h3d18;
mem_array[24487] = 16'h48da;
mem_array[24486] = 16'hbf81;
mem_array[24489] = 16'h48ce;
mem_array[24488] = 16'h3e61;
mem_array[24491] = 16'h1495;
mem_array[24490] = 16'h3cb1;
mem_array[24493] = 16'hcb9d;
mem_array[24492] = 16'hbe8b;
mem_array[24495] = 16'h2df1;
mem_array[24494] = 16'hbda0;
mem_array[24497] = 16'h550f;
mem_array[24496] = 16'h3d7f;
mem_array[24499] = 16'h10da;
mem_array[24498] = 16'h3e2d;
mem_array[24501] = 16'hcbbb;
mem_array[24500] = 16'hbda9;
mem_array[24503] = 16'h8b21;
mem_array[24502] = 16'h3ca2;
mem_array[24505] = 16'hfe3b;
mem_array[24504] = 16'hbea6;
mem_array[24507] = 16'hcc16;
mem_array[24506] = 16'h3ca9;
mem_array[24509] = 16'had42;
mem_array[24508] = 16'hbed6;
mem_array[24511] = 16'h9d8f;
mem_array[24510] = 16'h3e41;
mem_array[24513] = 16'h47ae;
mem_array[24512] = 16'h3b88;
mem_array[24515] = 16'h7c8d;
mem_array[24514] = 16'hbb80;
mem_array[24517] = 16'h39a9;
mem_array[24516] = 16'h3e92;
mem_array[24519] = 16'h9a9c;
mem_array[24518] = 16'hbd91;
mem_array[24521] = 16'hdb10;
mem_array[24520] = 16'h3e62;
mem_array[24523] = 16'h4dff;
mem_array[24522] = 16'h3e4f;
mem_array[24525] = 16'h7801;
mem_array[24524] = 16'h3da1;
mem_array[24527] = 16'ha69a;
mem_array[24526] = 16'h3d85;
mem_array[24529] = 16'h4364;
mem_array[24528] = 16'h3e72;
mem_array[24531] = 16'hbb8a;
mem_array[24530] = 16'hbe16;
mem_array[24533] = 16'h70ad;
mem_array[24532] = 16'h3d54;
mem_array[24535] = 16'h891b;
mem_array[24534] = 16'hbe26;
mem_array[24537] = 16'h1c59;
mem_array[24536] = 16'h3f1a;
mem_array[24539] = 16'h70bf;
mem_array[24538] = 16'h3e08;
mem_array[24541] = 16'h1829;
mem_array[24540] = 16'hbebd;
mem_array[24543] = 16'hcfc1;
mem_array[24542] = 16'h3d22;
mem_array[24545] = 16'hbe01;
mem_array[24544] = 16'hbbed;
mem_array[24547] = 16'h819d;
mem_array[24546] = 16'hbed5;
mem_array[24549] = 16'h4aa2;
mem_array[24548] = 16'h3d96;
mem_array[24551] = 16'hee9c;
mem_array[24550] = 16'hbeab;
mem_array[24553] = 16'he2c0;
mem_array[24552] = 16'hbe85;
mem_array[24555] = 16'h7a5f;
mem_array[24554] = 16'h3e07;
mem_array[24557] = 16'hd3f7;
mem_array[24556] = 16'hbc8d;
mem_array[24559] = 16'h4bc2;
mem_array[24558] = 16'hbeb1;
mem_array[24561] = 16'h4600;
mem_array[24560] = 16'hbde6;
mem_array[24563] = 16'h391b;
mem_array[24562] = 16'hbc5b;
mem_array[24565] = 16'h7cda;
mem_array[24564] = 16'hbddb;
mem_array[24567] = 16'hcf25;
mem_array[24566] = 16'h3cd8;
mem_array[24569] = 16'hd215;
mem_array[24568] = 16'hbea9;
mem_array[24571] = 16'h28e1;
mem_array[24570] = 16'h3ebf;
mem_array[24573] = 16'hf0b0;
mem_array[24572] = 16'hbe69;
mem_array[24575] = 16'h1204;
mem_array[24574] = 16'h3ec4;
mem_array[24577] = 16'h9285;
mem_array[24576] = 16'h3f00;
mem_array[24579] = 16'h329c;
mem_array[24578] = 16'h3ec6;
mem_array[24581] = 16'h00e3;
mem_array[24580] = 16'h3df6;
mem_array[24583] = 16'hda13;
mem_array[24582] = 16'h3f02;
mem_array[24585] = 16'h7e9b;
mem_array[24584] = 16'hbd90;
mem_array[24587] = 16'h39d3;
mem_array[24586] = 16'h3d2b;
mem_array[24589] = 16'h5508;
mem_array[24588] = 16'hbd8e;
mem_array[24591] = 16'h15e2;
mem_array[24590] = 16'hbbd5;
mem_array[24593] = 16'h59b6;
mem_array[24592] = 16'h3dab;
mem_array[24595] = 16'h4726;
mem_array[24594] = 16'hbdba;
mem_array[24597] = 16'hd3a5;
mem_array[24596] = 16'h3dd3;
mem_array[24599] = 16'h05e8;
mem_array[24598] = 16'h3e98;
mem_array[24601] = 16'hf22b;
mem_array[24600] = 16'hbee9;
mem_array[24603] = 16'h7c91;
mem_array[24602] = 16'hbb12;
mem_array[24605] = 16'h2e78;
mem_array[24604] = 16'h3e2f;
mem_array[24607] = 16'ha061;
mem_array[24606] = 16'hbe25;
mem_array[24609] = 16'h2614;
mem_array[24608] = 16'h3e96;
mem_array[24611] = 16'h0d64;
mem_array[24610] = 16'h3e05;
mem_array[24613] = 16'h0484;
mem_array[24612] = 16'hbe2b;
mem_array[24615] = 16'h428b;
mem_array[24614] = 16'hbe0a;
mem_array[24617] = 16'h4965;
mem_array[24616] = 16'h3da9;
mem_array[24619] = 16'h3a78;
mem_array[24618] = 16'hbf0a;
mem_array[24621] = 16'h2f38;
mem_array[24620] = 16'hbd72;
mem_array[24623] = 16'hf71f;
mem_array[24622] = 16'h3b39;
mem_array[24625] = 16'h0296;
mem_array[24624] = 16'hbe22;
mem_array[24627] = 16'h648f;
mem_array[24626] = 16'hbbba;
mem_array[24629] = 16'h4e5b;
mem_array[24628] = 16'hbdf5;
mem_array[24631] = 16'h446b;
mem_array[24630] = 16'h3e11;
mem_array[24633] = 16'h8680;
mem_array[24632] = 16'h3e4e;
mem_array[24635] = 16'h59fd;
mem_array[24634] = 16'h3e6b;
mem_array[24637] = 16'h4279;
mem_array[24636] = 16'h3e3b;
mem_array[24639] = 16'hfebe;
mem_array[24638] = 16'hbdaf;
mem_array[24641] = 16'hdbce;
mem_array[24640] = 16'h3dac;
mem_array[24643] = 16'h3bd9;
mem_array[24642] = 16'h3dc8;
mem_array[24645] = 16'hdf4f;
mem_array[24644] = 16'hbe87;
mem_array[24647] = 16'h0078;
mem_array[24646] = 16'h3e16;
mem_array[24649] = 16'he9b0;
mem_array[24648] = 16'h3d98;
mem_array[24651] = 16'hd802;
mem_array[24650] = 16'hbe67;
mem_array[24653] = 16'h4303;
mem_array[24652] = 16'hbe87;
mem_array[24655] = 16'h6c3b;
mem_array[24654] = 16'hbef3;
mem_array[24657] = 16'h15fc;
mem_array[24656] = 16'hbe4b;
mem_array[24659] = 16'h37f1;
mem_array[24658] = 16'h3d52;
mem_array[24661] = 16'h7f67;
mem_array[24660] = 16'hbe8e;
mem_array[24663] = 16'h9ef3;
mem_array[24662] = 16'h3e85;
mem_array[24665] = 16'hb35c;
mem_array[24664] = 16'h3d05;
mem_array[24667] = 16'h6063;
mem_array[24666] = 16'hbe90;
mem_array[24669] = 16'h6afa;
mem_array[24668] = 16'h3edf;
mem_array[24671] = 16'h61d5;
mem_array[24670] = 16'h3cc5;
mem_array[24673] = 16'h6c2a;
mem_array[24672] = 16'h3c57;
mem_array[24675] = 16'hb966;
mem_array[24674] = 16'h3982;
mem_array[24677] = 16'h4145;
mem_array[24676] = 16'hbc5a;
mem_array[24679] = 16'h0243;
mem_array[24678] = 16'h3efa;
mem_array[24681] = 16'heccd;
mem_array[24680] = 16'hbc82;
mem_array[24683] = 16'h92dd;
mem_array[24682] = 16'h3da6;
mem_array[24685] = 16'hd709;
mem_array[24684] = 16'h3d80;
mem_array[24687] = 16'h97fa;
mem_array[24686] = 16'hbe43;
mem_array[24689] = 16'he2a7;
mem_array[24688] = 16'hbda5;
mem_array[24691] = 16'h8870;
mem_array[24690] = 16'h3c98;
mem_array[24693] = 16'h73e2;
mem_array[24692] = 16'hbf53;
mem_array[24695] = 16'h5dca;
mem_array[24694] = 16'h3f0e;
mem_array[24697] = 16'h628e;
mem_array[24696] = 16'h3f01;
mem_array[24699] = 16'h58cd;
mem_array[24698] = 16'h3e43;
mem_array[24701] = 16'h0221;
mem_array[24700] = 16'h3ea1;
mem_array[24703] = 16'h84cb;
mem_array[24702] = 16'hbd8b;
mem_array[24705] = 16'hbb76;
mem_array[24704] = 16'h3e4f;
mem_array[24707] = 16'h3dac;
mem_array[24706] = 16'hbe8c;
mem_array[24709] = 16'h0c43;
mem_array[24708] = 16'hbd80;
mem_array[24711] = 16'h7bfb;
mem_array[24710] = 16'h3e3d;
mem_array[24713] = 16'he933;
mem_array[24712] = 16'hbed2;
mem_array[24715] = 16'h776d;
mem_array[24714] = 16'hbf70;
mem_array[24717] = 16'h8414;
mem_array[24716] = 16'hbe83;
mem_array[24719] = 16'h6159;
mem_array[24718] = 16'h3e26;
mem_array[24721] = 16'h1181;
mem_array[24720] = 16'hbea6;
mem_array[24723] = 16'h25a5;
mem_array[24722] = 16'hbe43;
mem_array[24725] = 16'hcc1c;
mem_array[24724] = 16'hbe1a;
mem_array[24727] = 16'h6a6c;
mem_array[24726] = 16'hbda6;
mem_array[24729] = 16'h34ff;
mem_array[24728] = 16'h3e2c;
mem_array[24731] = 16'h73ad;
mem_array[24730] = 16'hbe1a;
mem_array[24733] = 16'h16a9;
mem_array[24732] = 16'hbddf;
mem_array[24735] = 16'he44c;
mem_array[24734] = 16'hbc28;
mem_array[24737] = 16'he23f;
mem_array[24736] = 16'h3d2b;
mem_array[24739] = 16'h3f61;
mem_array[24738] = 16'h3d9e;
mem_array[24741] = 16'hde83;
mem_array[24740] = 16'h3c41;
mem_array[24743] = 16'hbaaa;
mem_array[24742] = 16'hba8f;
mem_array[24745] = 16'h161f;
mem_array[24744] = 16'h3ebe;
mem_array[24747] = 16'h58b6;
mem_array[24746] = 16'hbe92;
mem_array[24749] = 16'hf5af;
mem_array[24748] = 16'hbda8;
mem_array[24751] = 16'h4c54;
mem_array[24750] = 16'h3e1c;
mem_array[24753] = 16'h4092;
mem_array[24752] = 16'hbffc;
mem_array[24755] = 16'ha583;
mem_array[24754] = 16'h3e23;
mem_array[24757] = 16'hc9ed;
mem_array[24756] = 16'h3e83;
mem_array[24759] = 16'hb84d;
mem_array[24758] = 16'hbd7c;
mem_array[24761] = 16'h3557;
mem_array[24760] = 16'h3ecc;
mem_array[24763] = 16'h9344;
mem_array[24762] = 16'h3e91;
mem_array[24765] = 16'h98e5;
mem_array[24764] = 16'h3ee3;
mem_array[24767] = 16'h519c;
mem_array[24766] = 16'hbdcb;
mem_array[24769] = 16'hda24;
mem_array[24768] = 16'hbd98;
mem_array[24771] = 16'h2b52;
mem_array[24770] = 16'hbf3c;
mem_array[24773] = 16'h7fee;
mem_array[24772] = 16'h3e32;
mem_array[24775] = 16'hcc48;
mem_array[24774] = 16'hbfe1;
mem_array[24777] = 16'hb0a4;
mem_array[24776] = 16'hbdc2;
mem_array[24779] = 16'h5cc5;
mem_array[24778] = 16'h3ded;
mem_array[24781] = 16'hb5f3;
mem_array[24780] = 16'hbdba;
mem_array[24783] = 16'h99ae;
mem_array[24782] = 16'h3e08;
mem_array[24785] = 16'he833;
mem_array[24784] = 16'h3e06;
mem_array[24787] = 16'h51bb;
mem_array[24786] = 16'h3e21;
mem_array[24789] = 16'h1382;
mem_array[24788] = 16'hbd65;
mem_array[24791] = 16'hd180;
mem_array[24790] = 16'hbd1b;
mem_array[24793] = 16'h8058;
mem_array[24792] = 16'hbde9;
mem_array[24795] = 16'h0fed;
mem_array[24794] = 16'hbe31;
mem_array[24797] = 16'h8887;
mem_array[24796] = 16'hbe8a;
mem_array[24799] = 16'h929c;
mem_array[24798] = 16'hbf0b;
mem_array[24801] = 16'he26b;
mem_array[24800] = 16'h3d04;
mem_array[24803] = 16'h09a6;
mem_array[24802] = 16'hbd19;
mem_array[24805] = 16'h70fe;
mem_array[24804] = 16'h3e99;
mem_array[24807] = 16'hb74e;
mem_array[24806] = 16'hbe9c;
mem_array[24809] = 16'h66fb;
mem_array[24808] = 16'hbe86;
mem_array[24811] = 16'h5684;
mem_array[24810] = 16'hbc3e;
mem_array[24813] = 16'h487e;
mem_array[24812] = 16'hbfb8;
mem_array[24815] = 16'h078e;
mem_array[24814] = 16'h3e93;
mem_array[24817] = 16'haa54;
mem_array[24816] = 16'h3e71;
mem_array[24819] = 16'h9ae2;
mem_array[24818] = 16'hbd60;
mem_array[24821] = 16'hbb0f;
mem_array[24820] = 16'hbc96;
mem_array[24823] = 16'hdd38;
mem_array[24822] = 16'h3e94;
mem_array[24825] = 16'h9768;
mem_array[24824] = 16'h3e9e;
mem_array[24827] = 16'heb0c;
mem_array[24826] = 16'hbdb0;
mem_array[24829] = 16'h2cc4;
mem_array[24828] = 16'h3f14;
mem_array[24831] = 16'h795a;
mem_array[24830] = 16'hbdcb;
mem_array[24833] = 16'h9a5b;
mem_array[24832] = 16'hbced;
mem_array[24835] = 16'h34c4;
mem_array[24834] = 16'hc01a;
mem_array[24837] = 16'h79e6;
mem_array[24836] = 16'h3db8;
mem_array[24839] = 16'ha5e8;
mem_array[24838] = 16'hbe12;
mem_array[24841] = 16'hc86a;
mem_array[24840] = 16'h3eb2;
mem_array[24843] = 16'h803c;
mem_array[24842] = 16'hbde5;
mem_array[24845] = 16'hc934;
mem_array[24844] = 16'h3ddb;
mem_array[24847] = 16'h3930;
mem_array[24846] = 16'h3e91;
mem_array[24849] = 16'h86f1;
mem_array[24848] = 16'h3f05;
mem_array[24851] = 16'h640d;
mem_array[24850] = 16'h3e97;
mem_array[24853] = 16'ha5c1;
mem_array[24852] = 16'h3d80;
mem_array[24855] = 16'h7059;
mem_array[24854] = 16'hbbd1;
mem_array[24857] = 16'h5f48;
mem_array[24856] = 16'hbd42;
mem_array[24859] = 16'he2c0;
mem_array[24858] = 16'hbef6;
mem_array[24861] = 16'hc098;
mem_array[24860] = 16'hbd21;
mem_array[24863] = 16'h77ed;
mem_array[24862] = 16'h3d0c;
mem_array[24865] = 16'ha571;
mem_array[24864] = 16'h3ebd;
mem_array[24867] = 16'h293b;
mem_array[24866] = 16'h3de8;
mem_array[24869] = 16'h8b8e;
mem_array[24868] = 16'hbe88;
mem_array[24871] = 16'hfc2f;
mem_array[24870] = 16'h3d09;
mem_array[24873] = 16'hf138;
mem_array[24872] = 16'hbf76;
mem_array[24875] = 16'h9202;
mem_array[24874] = 16'h3e6c;
mem_array[24877] = 16'h4821;
mem_array[24876] = 16'h3d4e;
mem_array[24879] = 16'hc699;
mem_array[24878] = 16'hbe88;
mem_array[24881] = 16'hf2e2;
mem_array[24880] = 16'h3e6d;
mem_array[24883] = 16'h1f71;
mem_array[24882] = 16'h3cf6;
mem_array[24885] = 16'h2767;
mem_array[24884] = 16'h3f65;
mem_array[24887] = 16'haa8b;
mem_array[24886] = 16'h3e89;
mem_array[24889] = 16'h9b4b;
mem_array[24888] = 16'h3eb4;
mem_array[24891] = 16'hed41;
mem_array[24890] = 16'hbe1b;
mem_array[24893] = 16'hca5b;
mem_array[24892] = 16'hbee8;
mem_array[24895] = 16'h47ab;
mem_array[24894] = 16'hbfdb;
mem_array[24897] = 16'h387c;
mem_array[24896] = 16'hbc46;
mem_array[24899] = 16'h0010;
mem_array[24898] = 16'h3ead;
mem_array[24901] = 16'h821b;
mem_array[24900] = 16'hbe61;
mem_array[24903] = 16'h119f;
mem_array[24902] = 16'h3f23;
mem_array[24905] = 16'ha941;
mem_array[24904] = 16'hbe40;
mem_array[24907] = 16'h08f6;
mem_array[24906] = 16'h3e64;
mem_array[24909] = 16'hc2aa;
mem_array[24908] = 16'h3e1c;
mem_array[24911] = 16'h542c;
mem_array[24910] = 16'hbecb;
mem_array[24913] = 16'had15;
mem_array[24912] = 16'h3e58;
mem_array[24915] = 16'he505;
mem_array[24914] = 16'h3e89;
mem_array[24917] = 16'hdd48;
mem_array[24916] = 16'hbd48;
mem_array[24919] = 16'hedf0;
mem_array[24918] = 16'hbeda;
mem_array[24921] = 16'h3b64;
mem_array[24920] = 16'hbd8a;
mem_array[24923] = 16'h839e;
mem_array[24922] = 16'hbd5b;
mem_array[24925] = 16'h70b1;
mem_array[24924] = 16'h3ed9;
mem_array[24927] = 16'he7cd;
mem_array[24926] = 16'hbca3;
mem_array[24929] = 16'h92f4;
mem_array[24928] = 16'hbddf;
mem_array[24931] = 16'hece8;
mem_array[24930] = 16'hbd8b;
mem_array[24933] = 16'h00a1;
mem_array[24932] = 16'hbf60;
mem_array[24935] = 16'h854c;
mem_array[24934] = 16'hbe3a;
mem_array[24937] = 16'h9c07;
mem_array[24936] = 16'hbc6e;
mem_array[24939] = 16'h19b6;
mem_array[24938] = 16'hbe39;
mem_array[24941] = 16'h07f4;
mem_array[24940] = 16'h3e24;
mem_array[24943] = 16'h9541;
mem_array[24942] = 16'h3e7f;
mem_array[24945] = 16'h45f7;
mem_array[24944] = 16'h3d05;
mem_array[24947] = 16'h04ca;
mem_array[24946] = 16'h3eb9;
mem_array[24949] = 16'h8622;
mem_array[24948] = 16'h3e6d;
mem_array[24951] = 16'hee09;
mem_array[24950] = 16'h3ece;
mem_array[24953] = 16'hedc9;
mem_array[24952] = 16'hbe7b;
mem_array[24955] = 16'hc1bd;
mem_array[24954] = 16'hc013;
mem_array[24957] = 16'hdc88;
mem_array[24956] = 16'h3d22;
mem_array[24959] = 16'h9c3c;
mem_array[24958] = 16'hbe13;
mem_array[24961] = 16'he2d9;
mem_array[24960] = 16'h3f62;
mem_array[24963] = 16'h846d;
mem_array[24962] = 16'h3f13;
mem_array[24965] = 16'hfbea;
mem_array[24964] = 16'hbe9a;
mem_array[24967] = 16'ha06c;
mem_array[24966] = 16'h3f05;
mem_array[24969] = 16'h6521;
mem_array[24968] = 16'hbee6;
mem_array[24971] = 16'h0de0;
mem_array[24970] = 16'hbe56;
mem_array[24973] = 16'ha9c1;
mem_array[24972] = 16'h3f4d;
mem_array[24975] = 16'h078b;
mem_array[24974] = 16'hbf0a;
mem_array[24977] = 16'he7c6;
mem_array[24976] = 16'h3d83;
mem_array[24979] = 16'h9fb5;
mem_array[24978] = 16'hbede;
mem_array[24981] = 16'h6a6c;
mem_array[24980] = 16'h3d6e;
mem_array[24983] = 16'h34c5;
mem_array[24982] = 16'h3bf0;
mem_array[24985] = 16'hf4f8;
mem_array[24984] = 16'h3f08;
mem_array[24987] = 16'h645e;
mem_array[24986] = 16'h3e1a;
mem_array[24989] = 16'h3aa5;
mem_array[24988] = 16'h3e25;
mem_array[24991] = 16'h3b16;
mem_array[24990] = 16'h3eb1;
mem_array[24993] = 16'h6a3b;
mem_array[24992] = 16'hbed7;
mem_array[24995] = 16'h03fc;
mem_array[24994] = 16'hbe23;
mem_array[24997] = 16'h2dd6;
mem_array[24996] = 16'hbf29;
mem_array[24999] = 16'hf3f6;
mem_array[24998] = 16'hbece;
mem_array[25001] = 16'hf4db;
mem_array[25000] = 16'hbf22;
mem_array[25003] = 16'hb161;
mem_array[25002] = 16'h3d1c;
mem_array[25005] = 16'h4e06;
mem_array[25004] = 16'hbf84;
mem_array[25007] = 16'hc2cb;
mem_array[25006] = 16'h3f0e;
mem_array[25009] = 16'hd72c;
mem_array[25008] = 16'h3f45;
mem_array[25011] = 16'h68ba;
mem_array[25010] = 16'hbed6;
mem_array[25013] = 16'h27f0;
mem_array[25012] = 16'hbee6;
mem_array[25015] = 16'hedaa;
mem_array[25014] = 16'hbf43;
mem_array[25017] = 16'h42d4;
mem_array[25016] = 16'h3e0d;
mem_array[25019] = 16'h4796;
mem_array[25018] = 16'hbeba;
mem_array[25021] = 16'hb6fe;
mem_array[25020] = 16'h3f6a;
mem_array[25023] = 16'h1010;
mem_array[25022] = 16'h3f21;
mem_array[25025] = 16'hdb79;
mem_array[25024] = 16'h3d7a;
mem_array[25027] = 16'h1421;
mem_array[25026] = 16'h3ec0;
mem_array[25029] = 16'h9005;
mem_array[25028] = 16'h3f93;
mem_array[25031] = 16'h9f4a;
mem_array[25030] = 16'hbed5;
mem_array[25033] = 16'h274b;
mem_array[25032] = 16'h3f9c;
mem_array[25035] = 16'hbc0c;
mem_array[25034] = 16'hbd29;
mem_array[25037] = 16'h930e;
mem_array[25036] = 16'h3f02;
mem_array[25039] = 16'h251d;
mem_array[25038] = 16'h3e33;
mem_array[25041] = 16'h0bce;
mem_array[25040] = 16'hbcf6;
mem_array[25043] = 16'h3aa5;
mem_array[25042] = 16'h3c99;
mem_array[25045] = 16'h0b67;
mem_array[25044] = 16'h3ea2;
mem_array[25047] = 16'h3b4a;
mem_array[25046] = 16'hbccb;
mem_array[25049] = 16'hf656;
mem_array[25048] = 16'hbe93;
mem_array[25051] = 16'h6e3b;
mem_array[25050] = 16'h3ec0;
mem_array[25053] = 16'h0556;
mem_array[25052] = 16'hbe6b;
mem_array[25055] = 16'h2b07;
mem_array[25054] = 16'h3e2b;
mem_array[25057] = 16'h75aa;
mem_array[25056] = 16'h3eb7;
mem_array[25059] = 16'hefa7;
mem_array[25058] = 16'h3f14;
mem_array[25061] = 16'h3fe2;
mem_array[25060] = 16'h3e30;
mem_array[25063] = 16'ha22b;
mem_array[25062] = 16'hbefb;
mem_array[25065] = 16'h720e;
mem_array[25064] = 16'hbf40;
mem_array[25067] = 16'h20d2;
mem_array[25066] = 16'h3e1a;
mem_array[25069] = 16'h87b1;
mem_array[25068] = 16'h3edc;
mem_array[25071] = 16'hf1f6;
mem_array[25070] = 16'h3ee6;
mem_array[25073] = 16'hf382;
mem_array[25072] = 16'hbf0c;
mem_array[25075] = 16'hf370;
mem_array[25074] = 16'hbc95;
mem_array[25077] = 16'h7713;
mem_array[25076] = 16'h3ac0;
mem_array[25079] = 16'h6f7f;
mem_array[25078] = 16'hbec4;
mem_array[25081] = 16'h1c35;
mem_array[25080] = 16'hbf2e;
mem_array[25083] = 16'h3be1;
mem_array[25082] = 16'h3d63;
mem_array[25085] = 16'h9598;
mem_array[25084] = 16'h3f4f;
mem_array[25087] = 16'he0ed;
mem_array[25086] = 16'hbef0;
mem_array[25089] = 16'hcd85;
mem_array[25088] = 16'h3ef2;
mem_array[25091] = 16'h67c7;
mem_array[25090] = 16'hbe98;
mem_array[25093] = 16'h4612;
mem_array[25092] = 16'h3f80;
mem_array[25095] = 16'h87ea;
mem_array[25094] = 16'h3ef7;
mem_array[25097] = 16'h13e4;
mem_array[25096] = 16'h3f90;
mem_array[25099] = 16'h1852;
mem_array[25098] = 16'h3faf;
mem_array[25101] = 16'he70c;
mem_array[25100] = 16'hbdad;
mem_array[25103] = 16'h72d6;
mem_array[25102] = 16'h3d65;
mem_array[25105] = 16'ha786;
mem_array[25104] = 16'h3e8b;
mem_array[25107] = 16'h9e3e;
mem_array[25106] = 16'h3f2d;
mem_array[25109] = 16'h32b4;
mem_array[25108] = 16'h3e2e;
mem_array[25111] = 16'h00c5;
mem_array[25110] = 16'hbd32;
mem_array[25113] = 16'h13be;
mem_array[25112] = 16'h3f6c;
mem_array[25115] = 16'h5d65;
mem_array[25114] = 16'h3e43;
mem_array[25117] = 16'hb2ba;
mem_array[25116] = 16'hbf6e;
mem_array[25119] = 16'h7ee8;
mem_array[25118] = 16'h3ed3;
mem_array[25121] = 16'h1fbc;
mem_array[25120] = 16'hbf7e;
mem_array[25123] = 16'h9035;
mem_array[25122] = 16'hbf26;
mem_array[25125] = 16'h9e37;
mem_array[25124] = 16'hbeea;
mem_array[25127] = 16'h1651;
mem_array[25126] = 16'hbeaf;
mem_array[25129] = 16'h3f3c;
mem_array[25128] = 16'h3f61;
mem_array[25131] = 16'hdedb;
mem_array[25130] = 16'h3d01;
mem_array[25133] = 16'h747f;
mem_array[25132] = 16'h3efe;
mem_array[25135] = 16'h7a14;
mem_array[25134] = 16'hbdb0;
mem_array[25137] = 16'h1d26;
mem_array[25136] = 16'h3f39;
mem_array[25139] = 16'h24d5;
mem_array[25138] = 16'hbe21;
mem_array[25141] = 16'hf6ac;
mem_array[25140] = 16'h3c7a;
mem_array[25143] = 16'h144c;
mem_array[25142] = 16'hbd86;
mem_array[25145] = 16'h90f5;
mem_array[25144] = 16'h3ef2;
mem_array[25147] = 16'hf3d1;
mem_array[25146] = 16'hbcfb;
mem_array[25149] = 16'h6dea;
mem_array[25148] = 16'hbc83;
mem_array[25151] = 16'h082a;
mem_array[25150] = 16'hbda4;
mem_array[25153] = 16'h08a9;
mem_array[25152] = 16'h3ed0;
mem_array[25155] = 16'h1b45;
mem_array[25154] = 16'h3eac;
mem_array[25157] = 16'h5c7b;
mem_array[25156] = 16'h3f00;
mem_array[25159] = 16'hdf1e;
mem_array[25158] = 16'h3e70;
mem_array[25161] = 16'h8dd6;
mem_array[25160] = 16'h3dc0;
mem_array[25163] = 16'hc277;
mem_array[25162] = 16'hbcf4;
mem_array[25165] = 16'h61f3;
mem_array[25164] = 16'h3ca9;
mem_array[25167] = 16'h3b3e;
mem_array[25166] = 16'h3f06;
mem_array[25169] = 16'hb2c4;
mem_array[25168] = 16'h3de6;
mem_array[25171] = 16'h6f55;
mem_array[25170] = 16'hba40;
mem_array[25173] = 16'h8e06;
mem_array[25172] = 16'h3f0d;
mem_array[25175] = 16'h5806;
mem_array[25174] = 16'h3d24;
mem_array[25177] = 16'h05c8;
mem_array[25176] = 16'h3adb;
mem_array[25179] = 16'hc76d;
mem_array[25178] = 16'hbe22;
mem_array[25181] = 16'hc657;
mem_array[25180] = 16'hbe23;
mem_array[25183] = 16'h34b9;
mem_array[25182] = 16'hbe72;
mem_array[25185] = 16'h4477;
mem_array[25184] = 16'hbd19;
mem_array[25187] = 16'h2150;
mem_array[25186] = 16'hbece;
mem_array[25189] = 16'h057c;
mem_array[25188] = 16'h3ee8;
mem_array[25191] = 16'hf2e9;
mem_array[25190] = 16'h3ced;
mem_array[25193] = 16'h3c26;
mem_array[25192] = 16'h3ec3;
mem_array[25195] = 16'heca2;
mem_array[25194] = 16'hbd80;
mem_array[25197] = 16'h6189;
mem_array[25196] = 16'h3f0e;
mem_array[25199] = 16'hf6c1;
mem_array[25198] = 16'hbeb9;
mem_array[25201] = 16'hfd84;
mem_array[25200] = 16'hbc08;
mem_array[25203] = 16'hd7c5;
mem_array[25202] = 16'h3d0d;
mem_array[25205] = 16'ha2d4;
mem_array[25204] = 16'hbd1e;
mem_array[25207] = 16'hef82;
mem_array[25206] = 16'h3d1d;
mem_array[25209] = 16'h6a62;
mem_array[25208] = 16'hbdc9;
mem_array[25211] = 16'he339;
mem_array[25210] = 16'h3f20;
mem_array[25213] = 16'hd512;
mem_array[25212] = 16'h3e35;
mem_array[25215] = 16'hfd71;
mem_array[25214] = 16'h3e2d;
mem_array[25217] = 16'h05b1;
mem_array[25216] = 16'h3cbd;
mem_array[25219] = 16'hb383;
mem_array[25218] = 16'h3d40;
mem_array[25221] = 16'h0168;
mem_array[25220] = 16'h3d27;
mem_array[25223] = 16'h883e;
mem_array[25222] = 16'hbd44;
mem_array[25225] = 16'h3fef;
mem_array[25224] = 16'h3c9a;
mem_array[25227] = 16'h6f48;
mem_array[25226] = 16'h3d78;
mem_array[25229] = 16'he212;
mem_array[25228] = 16'hbd1b;
mem_array[25231] = 16'hd222;
mem_array[25230] = 16'hbea8;
mem_array[25233] = 16'hd708;
mem_array[25232] = 16'hbba2;
mem_array[25235] = 16'hece3;
mem_array[25234] = 16'h3d8b;
mem_array[25237] = 16'h2374;
mem_array[25236] = 16'hbe5c;
mem_array[25239] = 16'h6a57;
mem_array[25238] = 16'hbda0;
mem_array[25241] = 16'h54a8;
mem_array[25240] = 16'hbdbd;
mem_array[25243] = 16'h45d5;
mem_array[25242] = 16'h3f16;
mem_array[25245] = 16'hab20;
mem_array[25244] = 16'h3dc0;
mem_array[25247] = 16'h3f48;
mem_array[25246] = 16'h3dbb;
mem_array[25249] = 16'hf9be;
mem_array[25248] = 16'hbe06;
mem_array[25251] = 16'hb6af;
mem_array[25250] = 16'hbb97;
mem_array[25253] = 16'hb20d;
mem_array[25252] = 16'h3f67;
mem_array[25255] = 16'h1e10;
mem_array[25254] = 16'h3dc8;
mem_array[25257] = 16'h36cc;
mem_array[25256] = 16'h3dc3;
mem_array[25259] = 16'hbbce;
mem_array[25258] = 16'hbc88;
mem_array[25261] = 16'hda98;
mem_array[25260] = 16'h3d23;
mem_array[25263] = 16'h493c;
mem_array[25262] = 16'hbbf6;
mem_array[25265] = 16'h0e65;
mem_array[25264] = 16'hbd27;
mem_array[25267] = 16'h6050;
mem_array[25266] = 16'h3c8e;
mem_array[25269] = 16'h4866;
mem_array[25268] = 16'h3d12;
mem_array[25271] = 16'h5882;
mem_array[25270] = 16'h3d3e;
mem_array[25273] = 16'hdc28;
mem_array[25272] = 16'hbd1d;
mem_array[25275] = 16'h97bb;
mem_array[25274] = 16'hbbde;
mem_array[25277] = 16'h4625;
mem_array[25276] = 16'hbd06;
mem_array[25279] = 16'h4b09;
mem_array[25278] = 16'hbcf3;
mem_array[25281] = 16'h4847;
mem_array[25280] = 16'h3dc7;
mem_array[25283] = 16'h4f77;
mem_array[25282] = 16'hbd9f;
mem_array[25285] = 16'h2cf8;
mem_array[25284] = 16'h3d08;
mem_array[25287] = 16'h3e84;
mem_array[25286] = 16'hbe8c;
mem_array[25289] = 16'h0bfb;
mem_array[25288] = 16'hbd3a;
mem_array[25291] = 16'habd2;
mem_array[25290] = 16'hbe7a;
mem_array[25293] = 16'h39aa;
mem_array[25292] = 16'h3da5;
mem_array[25295] = 16'hc231;
mem_array[25294] = 16'h3d05;
mem_array[25297] = 16'hc0d1;
mem_array[25296] = 16'hbd49;
mem_array[25299] = 16'h3275;
mem_array[25298] = 16'h3d47;
mem_array[25301] = 16'haf3c;
mem_array[25300] = 16'h3c2e;
mem_array[25303] = 16'he5fe;
mem_array[25302] = 16'h3e98;
mem_array[25305] = 16'h1298;
mem_array[25304] = 16'h3d5c;
mem_array[25307] = 16'hc9dc;
mem_array[25306] = 16'hbcd7;
mem_array[25309] = 16'h7f3a;
mem_array[25308] = 16'h3e65;
mem_array[25311] = 16'h91d4;
mem_array[25310] = 16'hbd2c;
mem_array[25313] = 16'h1788;
mem_array[25312] = 16'h3dbc;
mem_array[25315] = 16'h6197;
mem_array[25314] = 16'hbda2;
mem_array[25317] = 16'hbf6a;
mem_array[25316] = 16'hbca8;
mem_array[25319] = 16'hf713;
mem_array[25318] = 16'h3d83;
mem_array[25321] = 16'hb48a;
mem_array[25320] = 16'h3ea4;
mem_array[25323] = 16'ha65a;
mem_array[25322] = 16'h3dd8;
mem_array[25325] = 16'h649f;
mem_array[25324] = 16'h3e52;
mem_array[25327] = 16'h5938;
mem_array[25326] = 16'hbdd4;
mem_array[25329] = 16'h9f8e;
mem_array[25328] = 16'hbca4;
mem_array[25331] = 16'h8b26;
mem_array[25330] = 16'hbde2;
mem_array[25333] = 16'hd5cd;
mem_array[25332] = 16'hbea3;
mem_array[25335] = 16'h7f07;
mem_array[25334] = 16'hbdb6;
mem_array[25337] = 16'hd7e2;
mem_array[25336] = 16'h3e16;
mem_array[25339] = 16'hd843;
mem_array[25338] = 16'hbda9;
mem_array[25341] = 16'h2f61;
mem_array[25340] = 16'h3b86;
mem_array[25343] = 16'h065b;
mem_array[25342] = 16'h3d9c;
mem_array[25345] = 16'h573f;
mem_array[25344] = 16'h3d1d;
mem_array[25347] = 16'h8629;
mem_array[25346] = 16'hbe8a;
mem_array[25349] = 16'h2fbe;
mem_array[25348] = 16'hbe73;
mem_array[25351] = 16'h95ef;
mem_array[25350] = 16'hbf15;
mem_array[25353] = 16'h854a;
mem_array[25352] = 16'h3f1d;
mem_array[25355] = 16'h1af4;
mem_array[25354] = 16'h3ef2;
mem_array[25357] = 16'haf18;
mem_array[25356] = 16'hbf73;
mem_array[25359] = 16'hd376;
mem_array[25358] = 16'h3f96;
mem_array[25361] = 16'h7fc4;
mem_array[25360] = 16'hbe21;
mem_array[25363] = 16'ha11b;
mem_array[25362] = 16'hbe91;
mem_array[25365] = 16'h0ade;
mem_array[25364] = 16'h3d58;
mem_array[25367] = 16'hd990;
mem_array[25366] = 16'hbe34;
mem_array[25369] = 16'hcf7a;
mem_array[25368] = 16'hbcca;
mem_array[25371] = 16'hf14f;
mem_array[25370] = 16'h3f35;
mem_array[25373] = 16'h1d7d;
mem_array[25372] = 16'h3e20;
mem_array[25375] = 16'h933c;
mem_array[25374] = 16'h3cc9;
mem_array[25377] = 16'hf7e9;
mem_array[25376] = 16'hbf19;
mem_array[25379] = 16'h89cf;
mem_array[25378] = 16'h3f95;
mem_array[25381] = 16'he53c;
mem_array[25380] = 16'h3e40;
mem_array[25383] = 16'h6efd;
mem_array[25382] = 16'h3f16;
mem_array[25385] = 16'h92ba;
mem_array[25384] = 16'hbef5;
mem_array[25387] = 16'h99d9;
mem_array[25386] = 16'hbf63;
mem_array[25389] = 16'he703;
mem_array[25388] = 16'h3f14;
mem_array[25391] = 16'h7266;
mem_array[25390] = 16'hbdb1;
mem_array[25393] = 16'hf26e;
mem_array[25392] = 16'h3e91;
mem_array[25395] = 16'hd8c4;
mem_array[25394] = 16'h3bd2;
mem_array[25397] = 16'h09d3;
mem_array[25396] = 16'hbec6;
mem_array[25399] = 16'h95ef;
mem_array[25398] = 16'hbe3a;
mem_array[25401] = 16'h9087;
mem_array[25400] = 16'hbd04;
mem_array[25403] = 16'h222c;
mem_array[25402] = 16'h3ca3;
mem_array[25405] = 16'h0075;
mem_array[25404] = 16'hbee2;
mem_array[25407] = 16'h1adc;
mem_array[25406] = 16'h3f35;
mem_array[25409] = 16'h6d2e;
mem_array[25408] = 16'hbe10;
mem_array[25411] = 16'h5c18;
mem_array[25410] = 16'h3f7d;
mem_array[25413] = 16'hf106;
mem_array[25412] = 16'h3df5;
mem_array[25415] = 16'h146e;
mem_array[25414] = 16'hbe3c;
mem_array[25417] = 16'h21ca;
mem_array[25416] = 16'hbda4;
mem_array[25419] = 16'h655e;
mem_array[25418] = 16'hbdfd;
mem_array[25421] = 16'hca12;
mem_array[25420] = 16'hbe55;
mem_array[25423] = 16'h74c6;
mem_array[25422] = 16'hbf66;
mem_array[25425] = 16'h47d3;
mem_array[25424] = 16'hbee3;
mem_array[25427] = 16'h2eea;
mem_array[25426] = 16'h3dae;
mem_array[25429] = 16'h2a44;
mem_array[25428] = 16'h3d2f;
mem_array[25431] = 16'h9502;
mem_array[25430] = 16'h3f8b;
mem_array[25433] = 16'hb7ca;
mem_array[25432] = 16'h3e8c;
mem_array[25435] = 16'h2a8a;
mem_array[25434] = 16'h3e7b;
mem_array[25437] = 16'h3b97;
mem_array[25436] = 16'h3da2;
mem_array[25439] = 16'h3866;
mem_array[25438] = 16'h3ed7;
mem_array[25441] = 16'hb24b;
mem_array[25440] = 16'h3ea4;
mem_array[25443] = 16'hdf39;
mem_array[25442] = 16'h3e54;
mem_array[25445] = 16'h270b;
mem_array[25444] = 16'h3c96;
mem_array[25447] = 16'hbdf2;
mem_array[25446] = 16'h3c0f;
mem_array[25449] = 16'h7c0b;
mem_array[25448] = 16'h3f15;
mem_array[25451] = 16'hc192;
mem_array[25450] = 16'hbf0e;
mem_array[25453] = 16'h4e27;
mem_array[25452] = 16'h3dd1;
mem_array[25455] = 16'hf6c6;
mem_array[25454] = 16'h3e06;
mem_array[25457] = 16'hec07;
mem_array[25456] = 16'hbedf;
mem_array[25459] = 16'h70ea;
mem_array[25458] = 16'h3f1f;
mem_array[25461] = 16'hdd5b;
mem_array[25460] = 16'hbcf6;
mem_array[25463] = 16'h83a4;
mem_array[25462] = 16'h3dc6;
mem_array[25465] = 16'h12ce;
mem_array[25464] = 16'h3df8;
mem_array[25467] = 16'hb64c;
mem_array[25466] = 16'h3f4e;
mem_array[25469] = 16'h967d;
mem_array[25468] = 16'hbe9d;
mem_array[25471] = 16'h9096;
mem_array[25470] = 16'h3ef6;
mem_array[25473] = 16'hdbef;
mem_array[25472] = 16'hbee4;
mem_array[25475] = 16'h3685;
mem_array[25474] = 16'h3f0e;
mem_array[25477] = 16'h58fb;
mem_array[25476] = 16'h3ee9;
mem_array[25479] = 16'h3a2c;
mem_array[25478] = 16'hbd77;
mem_array[25481] = 16'h48fc;
mem_array[25480] = 16'h3e7b;
mem_array[25483] = 16'hc809;
mem_array[25482] = 16'hbdb4;
mem_array[25485] = 16'h3bc5;
mem_array[25484] = 16'hbe2d;
mem_array[25487] = 16'hbbfe;
mem_array[25486] = 16'h3e3d;
mem_array[25489] = 16'hd3e3;
mem_array[25488] = 16'hbf20;
mem_array[25491] = 16'h8368;
mem_array[25490] = 16'h3ed8;
mem_array[25493] = 16'h7eb5;
mem_array[25492] = 16'hbef9;
mem_array[25495] = 16'h9f06;
mem_array[25494] = 16'h3e08;
mem_array[25497] = 16'hba8e;
mem_array[25496] = 16'h3f4c;
mem_array[25499] = 16'h60e2;
mem_array[25498] = 16'h3f04;
mem_array[25501] = 16'h1d45;
mem_array[25500] = 16'hbe8b;
mem_array[25503] = 16'h2ba2;
mem_array[25502] = 16'hbe59;
mem_array[25505] = 16'h134a;
mem_array[25504] = 16'hbec9;
mem_array[25507] = 16'h7a0f;
mem_array[25506] = 16'h3ed9;
mem_array[25509] = 16'hb633;
mem_array[25508] = 16'hbe02;
mem_array[25511] = 16'hef44;
mem_array[25510] = 16'hbf38;
mem_array[25513] = 16'h79ae;
mem_array[25512] = 16'hbee3;
mem_array[25515] = 16'h16f3;
mem_array[25514] = 16'h3eba;
mem_array[25517] = 16'h4270;
mem_array[25516] = 16'hbf8b;
mem_array[25519] = 16'ha42a;
mem_array[25518] = 16'hbeb1;
mem_array[25521] = 16'h670b;
mem_array[25520] = 16'hbcbd;
mem_array[25523] = 16'h010c;
mem_array[25522] = 16'h3dbd;
mem_array[25525] = 16'h3773;
mem_array[25524] = 16'h3e18;
mem_array[25527] = 16'hcbc2;
mem_array[25526] = 16'h3d35;
mem_array[25529] = 16'hf8ae;
mem_array[25528] = 16'hbf6d;
mem_array[25531] = 16'h6c18;
mem_array[25530] = 16'h3e13;
mem_array[25533] = 16'hb418;
mem_array[25532] = 16'hbef9;
mem_array[25535] = 16'h3944;
mem_array[25534] = 16'h3cea;
mem_array[25537] = 16'hacf7;
mem_array[25536] = 16'h3bfb;
mem_array[25539] = 16'hac43;
mem_array[25538] = 16'h3df1;
mem_array[25541] = 16'h0422;
mem_array[25540] = 16'h3def;
mem_array[25543] = 16'h0894;
mem_array[25542] = 16'h3e42;
mem_array[25545] = 16'he540;
mem_array[25544] = 16'hbe30;
mem_array[25547] = 16'hbccb;
mem_array[25546] = 16'h3e2d;
mem_array[25549] = 16'h1efd;
mem_array[25548] = 16'h3d15;
mem_array[25551] = 16'h438b;
mem_array[25550] = 16'h3f2f;
mem_array[25553] = 16'h66a4;
mem_array[25552] = 16'hbc2a;
mem_array[25555] = 16'h5106;
mem_array[25554] = 16'h3ede;
mem_array[25557] = 16'h78bc;
mem_array[25556] = 16'h3f59;
mem_array[25559] = 16'h2c63;
mem_array[25558] = 16'h3f3b;
mem_array[25561] = 16'hd7bf;
mem_array[25560] = 16'hbee7;
mem_array[25563] = 16'h408d;
mem_array[25562] = 16'h3ebd;
mem_array[25565] = 16'h08ab;
mem_array[25564] = 16'hbf74;
mem_array[25567] = 16'ha6ac;
mem_array[25566] = 16'h3ea8;
mem_array[25569] = 16'hd453;
mem_array[25568] = 16'hbc96;
mem_array[25571] = 16'h2412;
mem_array[25570] = 16'hbef5;
mem_array[25573] = 16'h1b0c;
mem_array[25572] = 16'h3d93;
mem_array[25575] = 16'heb88;
mem_array[25574] = 16'hbc14;
mem_array[25577] = 16'h925d;
mem_array[25576] = 16'hbf91;
mem_array[25579] = 16'hd3ae;
mem_array[25578] = 16'hbf57;
mem_array[25581] = 16'h26a7;
mem_array[25580] = 16'hbd88;
mem_array[25583] = 16'hd728;
mem_array[25582] = 16'h3c81;
mem_array[25585] = 16'h5f25;
mem_array[25584] = 16'h3e4b;
mem_array[25587] = 16'h845f;
mem_array[25586] = 16'h3f3f;
mem_array[25589] = 16'ha908;
mem_array[25588] = 16'hbe29;
mem_array[25591] = 16'h5668;
mem_array[25590] = 16'hbe43;
mem_array[25593] = 16'h31e3;
mem_array[25592] = 16'hbf66;
mem_array[25595] = 16'h8c3d;
mem_array[25594] = 16'h3e99;
mem_array[25597] = 16'h6763;
mem_array[25596] = 16'h3d7a;
mem_array[25599] = 16'h27bf;
mem_array[25598] = 16'h3e39;
mem_array[25601] = 16'h8b52;
mem_array[25600] = 16'hbe3e;
mem_array[25603] = 16'hf66a;
mem_array[25602] = 16'h3e6d;
mem_array[25605] = 16'h9f80;
mem_array[25604] = 16'h3ecf;
mem_array[25607] = 16'h2fc2;
mem_array[25606] = 16'h3e94;
mem_array[25609] = 16'h4d10;
mem_array[25608] = 16'hbbca;
mem_array[25611] = 16'h4847;
mem_array[25610] = 16'hbdde;
mem_array[25613] = 16'h74e4;
mem_array[25612] = 16'h3de5;
mem_array[25615] = 16'h2123;
mem_array[25614] = 16'h3ea6;
mem_array[25617] = 16'h8765;
mem_array[25616] = 16'h3edc;
mem_array[25619] = 16'h352c;
mem_array[25618] = 16'h3e62;
mem_array[25621] = 16'h4798;
mem_array[25620] = 16'hbcd8;
mem_array[25623] = 16'h9afe;
mem_array[25622] = 16'h3e45;
mem_array[25625] = 16'h426d;
mem_array[25624] = 16'hbfb0;
mem_array[25627] = 16'h9568;
mem_array[25626] = 16'h3f4b;
mem_array[25629] = 16'hd1b7;
mem_array[25628] = 16'h3e89;
mem_array[25631] = 16'h853b;
mem_array[25630] = 16'hbf3a;
mem_array[25633] = 16'h4418;
mem_array[25632] = 16'hbea8;
mem_array[25635] = 16'haa04;
mem_array[25634] = 16'hbe71;
mem_array[25637] = 16'h5cc7;
mem_array[25636] = 16'hbeff;
mem_array[25639] = 16'h79b9;
mem_array[25638] = 16'hbeb6;
mem_array[25641] = 16'hfc78;
mem_array[25640] = 16'hbd95;
mem_array[25643] = 16'h59d5;
mem_array[25642] = 16'hbdb1;
mem_array[25645] = 16'h684c;
mem_array[25644] = 16'h3eaf;
mem_array[25647] = 16'h98fb;
mem_array[25646] = 16'h3e08;
mem_array[25649] = 16'h427a;
mem_array[25648] = 16'hbf0f;
mem_array[25651] = 16'h04f0;
mem_array[25650] = 16'h3e12;
mem_array[25653] = 16'hfb81;
mem_array[25652] = 16'hbe07;
mem_array[25655] = 16'h8de6;
mem_array[25654] = 16'h3c64;
mem_array[25657] = 16'hfcb4;
mem_array[25656] = 16'hbe07;
mem_array[25659] = 16'h00cc;
mem_array[25658] = 16'hbe0c;
mem_array[25661] = 16'hdc40;
mem_array[25660] = 16'h3e3f;
mem_array[25663] = 16'h63a8;
mem_array[25662] = 16'h3d52;
mem_array[25665] = 16'hc8cb;
mem_array[25664] = 16'h3eed;
mem_array[25667] = 16'h26d9;
mem_array[25666] = 16'h3e99;
mem_array[25669] = 16'h1da9;
mem_array[25668] = 16'hbd84;
mem_array[25671] = 16'h1558;
mem_array[25670] = 16'hbc1b;
mem_array[25673] = 16'h09ae;
mem_array[25672] = 16'hbd7e;
mem_array[25675] = 16'hde89;
mem_array[25674] = 16'h3ba7;
mem_array[25677] = 16'h133d;
mem_array[25676] = 16'h3db7;
mem_array[25679] = 16'h3c29;
mem_array[25678] = 16'h3f04;
mem_array[25681] = 16'h5934;
mem_array[25680] = 16'h3e98;
mem_array[25683] = 16'he592;
mem_array[25682] = 16'hbcb1;
mem_array[25685] = 16'h560f;
mem_array[25684] = 16'hc028;
mem_array[25687] = 16'h30c8;
mem_array[25686] = 16'h3e86;
mem_array[25689] = 16'haef2;
mem_array[25688] = 16'hbdb9;
mem_array[25691] = 16'h3dd8;
mem_array[25690] = 16'hbf13;
mem_array[25693] = 16'h8b81;
mem_array[25692] = 16'hbf36;
mem_array[25695] = 16'haa75;
mem_array[25694] = 16'hbf12;
mem_array[25697] = 16'hef79;
mem_array[25696] = 16'hbe9f;
mem_array[25699] = 16'h8a12;
mem_array[25698] = 16'h3dcb;
mem_array[25701] = 16'h39bd;
mem_array[25700] = 16'hbdb0;
mem_array[25703] = 16'h684f;
mem_array[25702] = 16'h3d0d;
mem_array[25705] = 16'h3fa7;
mem_array[25704] = 16'h3ec3;
mem_array[25707] = 16'h4b6a;
mem_array[25706] = 16'h3ef7;
mem_array[25709] = 16'hc134;
mem_array[25708] = 16'hbe3f;
mem_array[25711] = 16'h9683;
mem_array[25710] = 16'hbdc7;
mem_array[25713] = 16'hdb3a;
mem_array[25712] = 16'h3e20;
mem_array[25715] = 16'hab30;
mem_array[25714] = 16'h3dc2;
mem_array[25717] = 16'h362f;
mem_array[25716] = 16'h3e5f;
mem_array[25719] = 16'hf1fe;
mem_array[25718] = 16'h3e65;
mem_array[25721] = 16'h87e4;
mem_array[25720] = 16'h3e63;
mem_array[25723] = 16'hd143;
mem_array[25722] = 16'h3ddd;
mem_array[25725] = 16'h6843;
mem_array[25724] = 16'h3ed4;
mem_array[25727] = 16'h2ae5;
mem_array[25726] = 16'h3e8a;
mem_array[25729] = 16'h52f1;
mem_array[25728] = 16'hbe14;
mem_array[25731] = 16'h04b2;
mem_array[25730] = 16'hbf32;
mem_array[25733] = 16'h4421;
mem_array[25732] = 16'hbe34;
mem_array[25735] = 16'h52cf;
mem_array[25734] = 16'h3e24;
mem_array[25737] = 16'hf332;
mem_array[25736] = 16'hbda4;
mem_array[25739] = 16'ha52b;
mem_array[25738] = 16'h3ef1;
mem_array[25741] = 16'hca2b;
mem_array[25740] = 16'h3e74;
mem_array[25743] = 16'h4bc1;
mem_array[25742] = 16'h3e89;
mem_array[25745] = 16'hff70;
mem_array[25744] = 16'hbfbb;
mem_array[25747] = 16'hc8b6;
mem_array[25746] = 16'h3ebe;
mem_array[25749] = 16'haad7;
mem_array[25748] = 16'h3d84;
mem_array[25751] = 16'h141d;
mem_array[25750] = 16'hbe27;
mem_array[25753] = 16'h263f;
mem_array[25752] = 16'hbeff;
mem_array[25755] = 16'hc292;
mem_array[25754] = 16'hbe9c;
mem_array[25757] = 16'h2dcc;
mem_array[25756] = 16'hbcdf;
mem_array[25759] = 16'h1c6d;
mem_array[25758] = 16'h3f1a;
mem_array[25761] = 16'h0827;
mem_array[25760] = 16'hbe0a;
mem_array[25763] = 16'hb9fd;
mem_array[25762] = 16'h3da1;
mem_array[25765] = 16'h4649;
mem_array[25764] = 16'h3e95;
mem_array[25767] = 16'h3135;
mem_array[25766] = 16'h3f48;
mem_array[25769] = 16'h20c4;
mem_array[25768] = 16'h3e23;
mem_array[25771] = 16'hc73a;
mem_array[25770] = 16'hbc05;
mem_array[25773] = 16'h5b93;
mem_array[25772] = 16'h3f04;
mem_array[25775] = 16'hf154;
mem_array[25774] = 16'h3b47;
mem_array[25777] = 16'h330e;
mem_array[25776] = 16'h3ca3;
mem_array[25779] = 16'h965b;
mem_array[25778] = 16'h3e06;
mem_array[25781] = 16'h8831;
mem_array[25780] = 16'hbd26;
mem_array[25783] = 16'h9a2b;
mem_array[25782] = 16'hbd31;
mem_array[25785] = 16'hc4cb;
mem_array[25784] = 16'h3eee;
mem_array[25787] = 16'hc2e2;
mem_array[25786] = 16'h3d73;
mem_array[25789] = 16'hf71c;
mem_array[25788] = 16'h3e51;
mem_array[25791] = 16'h20f9;
mem_array[25790] = 16'hbf61;
mem_array[25793] = 16'ha35c;
mem_array[25792] = 16'hbcdc;
mem_array[25795] = 16'hc384;
mem_array[25794] = 16'h3d9c;
mem_array[25797] = 16'h88e9;
mem_array[25796] = 16'hbe00;
mem_array[25799] = 16'h5102;
mem_array[25798] = 16'h3edd;
mem_array[25801] = 16'h79ca;
mem_array[25800] = 16'hbd67;
mem_array[25803] = 16'ha23c;
mem_array[25802] = 16'h3f29;
mem_array[25805] = 16'he6bc;
mem_array[25804] = 16'hbee4;
mem_array[25807] = 16'h6532;
mem_array[25806] = 16'h3e3a;
mem_array[25809] = 16'h9d66;
mem_array[25808] = 16'hbe50;
mem_array[25811] = 16'h1b8e;
mem_array[25810] = 16'hbd9a;
mem_array[25813] = 16'hf43d;
mem_array[25812] = 16'hbe6c;
mem_array[25815] = 16'h5167;
mem_array[25814] = 16'hbe86;
mem_array[25817] = 16'h76f8;
mem_array[25816] = 16'h3e00;
mem_array[25819] = 16'h740b;
mem_array[25818] = 16'hbf3c;
mem_array[25821] = 16'h4be7;
mem_array[25820] = 16'hbc4e;
mem_array[25823] = 16'h2041;
mem_array[25822] = 16'hbd8a;
mem_array[25825] = 16'h9ed3;
mem_array[25824] = 16'h3dfe;
mem_array[25827] = 16'ha52a;
mem_array[25826] = 16'h3e8c;
mem_array[25829] = 16'h1f8c;
mem_array[25828] = 16'h3e26;
mem_array[25831] = 16'h91cb;
mem_array[25830] = 16'h3d1d;
mem_array[25833] = 16'h6af4;
mem_array[25832] = 16'h3ecc;
mem_array[25835] = 16'hd7ef;
mem_array[25834] = 16'h3e7b;
mem_array[25837] = 16'h331b;
mem_array[25836] = 16'h3e11;
mem_array[25839] = 16'hc93c;
mem_array[25838] = 16'h3e81;
mem_array[25841] = 16'hc2e5;
mem_array[25840] = 16'hbd6a;
mem_array[25843] = 16'h9fc3;
mem_array[25842] = 16'hbd8f;
mem_array[25845] = 16'h801d;
mem_array[25844] = 16'h3ea6;
mem_array[25847] = 16'hc8b1;
mem_array[25846] = 16'h3dee;
mem_array[25849] = 16'hb52a;
mem_array[25848] = 16'h3e1f;
mem_array[25851] = 16'h2fab;
mem_array[25850] = 16'hbf35;
mem_array[25853] = 16'h58f5;
mem_array[25852] = 16'hbe70;
mem_array[25855] = 16'h8f6e;
mem_array[25854] = 16'h3e6f;
mem_array[25857] = 16'hffae;
mem_array[25856] = 16'h3d4a;
mem_array[25859] = 16'h2da2;
mem_array[25858] = 16'h3f2b;
mem_array[25861] = 16'hc3c9;
mem_array[25860] = 16'h3eac;
mem_array[25863] = 16'h9746;
mem_array[25862] = 16'h3e19;
mem_array[25865] = 16'h1ed9;
mem_array[25864] = 16'h3e1e;
mem_array[25867] = 16'hf91d;
mem_array[25866] = 16'h3e56;
mem_array[25869] = 16'hf5df;
mem_array[25868] = 16'hbdf6;
mem_array[25871] = 16'h3c5e;
mem_array[25870] = 16'hbeb8;
mem_array[25873] = 16'h538e;
mem_array[25872] = 16'hbe14;
mem_array[25875] = 16'hc08f;
mem_array[25874] = 16'hbee1;
mem_array[25877] = 16'h8cdc;
mem_array[25876] = 16'h3e09;
mem_array[25879] = 16'h4d49;
mem_array[25878] = 16'h3e70;
mem_array[25881] = 16'h8500;
mem_array[25880] = 16'hbc88;
mem_array[25883] = 16'h6e56;
mem_array[25882] = 16'h3d23;
mem_array[25885] = 16'he8ab;
mem_array[25884] = 16'h3eb1;
mem_array[25887] = 16'hc951;
mem_array[25886] = 16'h3dfc;
mem_array[25889] = 16'h0968;
mem_array[25888] = 16'h3f16;
mem_array[25891] = 16'h012f;
mem_array[25890] = 16'h3cbe;
mem_array[25893] = 16'h88e5;
mem_array[25892] = 16'h3dea;
mem_array[25895] = 16'h08d5;
mem_array[25894] = 16'hbccd;
mem_array[25897] = 16'hd3c5;
mem_array[25896] = 16'h3dc4;
mem_array[25899] = 16'h5e5c;
mem_array[25898] = 16'h3dda;
mem_array[25901] = 16'hf4ad;
mem_array[25900] = 16'h3dec;
mem_array[25903] = 16'h6b28;
mem_array[25902] = 16'hbdd0;
mem_array[25905] = 16'hd674;
mem_array[25904] = 16'h3d43;
mem_array[25907] = 16'hc904;
mem_array[25906] = 16'hbe03;
mem_array[25909] = 16'h425b;
mem_array[25908] = 16'h3e45;
mem_array[25911] = 16'h698a;
mem_array[25910] = 16'hbf2a;
mem_array[25913] = 16'h5d27;
mem_array[25912] = 16'h3d53;
mem_array[25915] = 16'h3efd;
mem_array[25914] = 16'h3bca;
mem_array[25917] = 16'h70bb;
mem_array[25916] = 16'h3caf;
mem_array[25919] = 16'hbfd4;
mem_array[25918] = 16'h3eb9;
mem_array[25921] = 16'had00;
mem_array[25920] = 16'h3e4e;
mem_array[25923] = 16'h1d4b;
mem_array[25922] = 16'hc010;
mem_array[25925] = 16'he736;
mem_array[25924] = 16'hbd40;
mem_array[25927] = 16'h1189;
mem_array[25926] = 16'hbe05;
mem_array[25929] = 16'h1bae;
mem_array[25928] = 16'hbdb2;
mem_array[25931] = 16'h4e62;
mem_array[25930] = 16'h3cbd;
mem_array[25933] = 16'hcafc;
mem_array[25932] = 16'h3d3d;
mem_array[25935] = 16'h2766;
mem_array[25934] = 16'hbeb6;
mem_array[25937] = 16'h96ed;
mem_array[25936] = 16'h3eb0;
mem_array[25939] = 16'hd428;
mem_array[25938] = 16'h3e16;
mem_array[25941] = 16'h73b6;
mem_array[25940] = 16'hbdc2;
mem_array[25943] = 16'heba3;
mem_array[25942] = 16'h3bb5;
mem_array[25945] = 16'hddfc;
mem_array[25944] = 16'h3cab;
mem_array[25947] = 16'hf454;
mem_array[25946] = 16'hb9f3;
mem_array[25949] = 16'hb5ad;
mem_array[25948] = 16'h3ed1;
mem_array[25951] = 16'hf6cb;
mem_array[25950] = 16'h3a94;
mem_array[25953] = 16'hf184;
mem_array[25952] = 16'hbdaf;
mem_array[25955] = 16'h992a;
mem_array[25954] = 16'hbe79;
mem_array[25957] = 16'ha592;
mem_array[25956] = 16'hbea9;
mem_array[25959] = 16'hac92;
mem_array[25958] = 16'h3e97;
mem_array[25961] = 16'h0216;
mem_array[25960] = 16'hbdff;
mem_array[25963] = 16'hd296;
mem_array[25962] = 16'hbe87;
mem_array[25965] = 16'hc5f1;
mem_array[25964] = 16'h3e78;
mem_array[25967] = 16'hafac;
mem_array[25966] = 16'h3c95;
mem_array[25969] = 16'hee08;
mem_array[25968] = 16'h3e94;
mem_array[25971] = 16'h4e9a;
mem_array[25970] = 16'hbf53;
mem_array[25973] = 16'h577d;
mem_array[25972] = 16'h3ca4;
mem_array[25975] = 16'hc80d;
mem_array[25974] = 16'hbe2c;
mem_array[25977] = 16'h530e;
mem_array[25976] = 16'hbe40;
mem_array[25979] = 16'h4e68;
mem_array[25978] = 16'h3cc4;
mem_array[25981] = 16'h7daa;
mem_array[25980] = 16'h3de7;
mem_array[25983] = 16'he717;
mem_array[25982] = 16'hbff4;
mem_array[25985] = 16'hdf31;
mem_array[25984] = 16'hbe68;
mem_array[25987] = 16'hdc4e;
mem_array[25986] = 16'hbf03;
mem_array[25989] = 16'h5d2e;
mem_array[25988] = 16'hbe21;
mem_array[25991] = 16'he4c4;
mem_array[25990] = 16'h3dd7;
mem_array[25993] = 16'h7810;
mem_array[25992] = 16'h3e75;
mem_array[25995] = 16'h4722;
mem_array[25994] = 16'hbeac;
mem_array[25997] = 16'h5892;
mem_array[25996] = 16'h3e94;
mem_array[25999] = 16'h783c;
mem_array[25998] = 16'h3e32;
mem_array[26001] = 16'h78bd;
mem_array[26000] = 16'hbb70;
mem_array[26003] = 16'hd5ad;
mem_array[26002] = 16'hbcad;
mem_array[26005] = 16'he219;
mem_array[26004] = 16'hbec9;
mem_array[26007] = 16'h02db;
mem_array[26006] = 16'h3d96;
mem_array[26009] = 16'hbc82;
mem_array[26008] = 16'h3e49;
mem_array[26011] = 16'hb158;
mem_array[26010] = 16'h3e61;
mem_array[26013] = 16'h22e7;
mem_array[26012] = 16'h3d9d;
mem_array[26015] = 16'hb308;
mem_array[26014] = 16'h3ac2;
mem_array[26017] = 16'h84dd;
mem_array[26016] = 16'hbe9c;
mem_array[26019] = 16'h702b;
mem_array[26018] = 16'h3c38;
mem_array[26021] = 16'hb324;
mem_array[26020] = 16'h3da8;
mem_array[26023] = 16'h4f19;
mem_array[26022] = 16'hbd31;
mem_array[26025] = 16'h7fc8;
mem_array[26024] = 16'hbdcd;
mem_array[26027] = 16'h2681;
mem_array[26026] = 16'hbd9b;
mem_array[26029] = 16'h3ee3;
mem_array[26028] = 16'h3e99;
mem_array[26031] = 16'hd2a4;
mem_array[26030] = 16'hbe3c;
mem_array[26033] = 16'he1e8;
mem_array[26032] = 16'h3e04;
mem_array[26035] = 16'h6cb9;
mem_array[26034] = 16'hbd86;
mem_array[26037] = 16'h34f3;
mem_array[26036] = 16'hbe75;
mem_array[26039] = 16'hc51a;
mem_array[26038] = 16'hbe0e;
mem_array[26041] = 16'h9acd;
mem_array[26040] = 16'hbe7b;
mem_array[26043] = 16'h594d;
mem_array[26042] = 16'hbf0b;
mem_array[26045] = 16'hebe1;
mem_array[26044] = 16'hbdb7;
mem_array[26047] = 16'h4d95;
mem_array[26046] = 16'hbf83;
mem_array[26049] = 16'h0d98;
mem_array[26048] = 16'h3e8b;
mem_array[26051] = 16'hd50e;
mem_array[26050] = 16'hbd0c;
mem_array[26053] = 16'h7d32;
mem_array[26052] = 16'h3ead;
mem_array[26055] = 16'hfe50;
mem_array[26054] = 16'hbe65;
mem_array[26057] = 16'h69a1;
mem_array[26056] = 16'h3cab;
mem_array[26059] = 16'h4d23;
mem_array[26058] = 16'h3d88;
mem_array[26061] = 16'h2663;
mem_array[26060] = 16'h3d97;
mem_array[26063] = 16'hc4b2;
mem_array[26062] = 16'hbca7;
mem_array[26065] = 16'hfb08;
mem_array[26064] = 16'hbdb9;
mem_array[26067] = 16'hc15b;
mem_array[26066] = 16'h3e1b;
mem_array[26069] = 16'h2b49;
mem_array[26068] = 16'h3c69;
mem_array[26071] = 16'he3a2;
mem_array[26070] = 16'h3eb1;
mem_array[26073] = 16'h3198;
mem_array[26072] = 16'hbe0e;
mem_array[26075] = 16'he3d7;
mem_array[26074] = 16'hbd8f;
mem_array[26077] = 16'h6e9c;
mem_array[26076] = 16'h3db5;
mem_array[26079] = 16'hafb9;
mem_array[26078] = 16'hbead;
mem_array[26081] = 16'ha08d;
mem_array[26080] = 16'h3e26;
mem_array[26083] = 16'ha463;
mem_array[26082] = 16'h3e5f;
mem_array[26085] = 16'h8b0f;
mem_array[26084] = 16'hbefd;
mem_array[26087] = 16'hdce5;
mem_array[26086] = 16'h3d9e;
mem_array[26089] = 16'h1026;
mem_array[26088] = 16'h3ca1;
mem_array[26091] = 16'h7350;
mem_array[26090] = 16'h3dcd;
mem_array[26093] = 16'h601b;
mem_array[26092] = 16'h3e5e;
mem_array[26095] = 16'h2d53;
mem_array[26094] = 16'hbdd3;
mem_array[26097] = 16'hbbe9;
mem_array[26096] = 16'hbe80;
mem_array[26099] = 16'hd227;
mem_array[26098] = 16'h3d3c;
mem_array[26101] = 16'h2338;
mem_array[26100] = 16'hbe55;
mem_array[26103] = 16'h5a83;
mem_array[26102] = 16'h3dc4;
mem_array[26105] = 16'h23a3;
mem_array[26104] = 16'hbc90;
mem_array[26107] = 16'h6dc6;
mem_array[26106] = 16'hbf7f;
mem_array[26109] = 16'h202b;
mem_array[26108] = 16'h3e6f;
mem_array[26111] = 16'he162;
mem_array[26110] = 16'hbd98;
mem_array[26113] = 16'h65af;
mem_array[26112] = 16'h3d52;
mem_array[26115] = 16'h72ba;
mem_array[26114] = 16'hbea7;
mem_array[26117] = 16'h628b;
mem_array[26116] = 16'hbc9f;
mem_array[26119] = 16'h9a40;
mem_array[26118] = 16'hbebc;
mem_array[26121] = 16'h031e;
mem_array[26120] = 16'hbc9b;
mem_array[26123] = 16'h872a;
mem_array[26122] = 16'h3d6d;
mem_array[26125] = 16'h1283;
mem_array[26124] = 16'hbe03;
mem_array[26127] = 16'h195d;
mem_array[26126] = 16'hbe7c;
mem_array[26129] = 16'had22;
mem_array[26128] = 16'hbe34;
mem_array[26131] = 16'he4dc;
mem_array[26130] = 16'h3e91;
mem_array[26133] = 16'hcab0;
mem_array[26132] = 16'hbe57;
mem_array[26135] = 16'hc4c2;
mem_array[26134] = 16'hbded;
mem_array[26137] = 16'h34b4;
mem_array[26136] = 16'h3e94;
mem_array[26139] = 16'hf1f3;
mem_array[26138] = 16'hbee8;
mem_array[26141] = 16'hf2ac;
mem_array[26140] = 16'h3f05;
mem_array[26143] = 16'hf1b8;
mem_array[26142] = 16'h3ea4;
mem_array[26145] = 16'h4094;
mem_array[26144] = 16'hbe4f;
mem_array[26147] = 16'h5889;
mem_array[26146] = 16'h3bca;
mem_array[26149] = 16'h3ac0;
mem_array[26148] = 16'h3dc8;
mem_array[26151] = 16'h3681;
mem_array[26150] = 16'hbbb6;
mem_array[26153] = 16'hfeac;
mem_array[26152] = 16'h3e0a;
mem_array[26155] = 16'h3cbb;
mem_array[26154] = 16'hbe18;
mem_array[26157] = 16'h8872;
mem_array[26156] = 16'h3d8d;
mem_array[26159] = 16'he305;
mem_array[26158] = 16'h3db6;
mem_array[26161] = 16'h4373;
mem_array[26160] = 16'h3da9;
mem_array[26163] = 16'h3413;
mem_array[26162] = 16'hbe26;
mem_array[26165] = 16'h2b91;
mem_array[26164] = 16'h3dca;
mem_array[26167] = 16'hd7a5;
mem_array[26166] = 16'hbeba;
mem_array[26169] = 16'ha6e5;
mem_array[26168] = 16'hbe79;
mem_array[26171] = 16'he40d;
mem_array[26170] = 16'hbdda;
mem_array[26173] = 16'h3fb8;
mem_array[26172] = 16'hbe96;
mem_array[26175] = 16'hd322;
mem_array[26174] = 16'hbe59;
mem_array[26177] = 16'he422;
mem_array[26176] = 16'h3ebc;
mem_array[26179] = 16'h02fd;
mem_array[26178] = 16'h3eb5;
mem_array[26181] = 16'hb9f7;
mem_array[26180] = 16'hbdbe;
mem_array[26183] = 16'h3660;
mem_array[26182] = 16'hbd33;
mem_array[26185] = 16'h6a07;
mem_array[26184] = 16'hbd64;
mem_array[26187] = 16'h84ac;
mem_array[26186] = 16'h3d4e;
mem_array[26189] = 16'h2346;
mem_array[26188] = 16'hba02;
mem_array[26191] = 16'h1554;
mem_array[26190] = 16'h3e05;
mem_array[26193] = 16'h5a7b;
mem_array[26192] = 16'h3eb0;
mem_array[26195] = 16'h8403;
mem_array[26194] = 16'h3ce6;
mem_array[26197] = 16'h00d2;
mem_array[26196] = 16'h3ebb;
mem_array[26199] = 16'h20ea;
mem_array[26198] = 16'h3ca0;
mem_array[26201] = 16'h3a7c;
mem_array[26200] = 16'h3e78;
mem_array[26203] = 16'h96d2;
mem_array[26202] = 16'hbd10;
mem_array[26205] = 16'h921c;
mem_array[26204] = 16'h3e44;
mem_array[26207] = 16'he42d;
mem_array[26206] = 16'hbd08;
mem_array[26209] = 16'h4ea6;
mem_array[26208] = 16'h3c58;
mem_array[26211] = 16'hf9a6;
mem_array[26210] = 16'hbda8;
mem_array[26213] = 16'h23ad;
mem_array[26212] = 16'hbcbb;
mem_array[26215] = 16'hc21b;
mem_array[26214] = 16'hbda8;
mem_array[26217] = 16'ha86c;
mem_array[26216] = 16'h3ee1;
mem_array[26219] = 16'h56ef;
mem_array[26218] = 16'h3e82;
mem_array[26221] = 16'ha48d;
mem_array[26220] = 16'hbd9a;
mem_array[26223] = 16'h6b67;
mem_array[26222] = 16'h3ddd;
mem_array[26225] = 16'ha0e8;
mem_array[26224] = 16'h3dfd;
mem_array[26227] = 16'h1f59;
mem_array[26226] = 16'hbf0f;
mem_array[26229] = 16'h1573;
mem_array[26228] = 16'h3e67;
mem_array[26231] = 16'h8751;
mem_array[26230] = 16'hbe8c;
mem_array[26233] = 16'hac7c;
mem_array[26232] = 16'hbd54;
mem_array[26235] = 16'h68c1;
mem_array[26234] = 16'h3dd5;
mem_array[26237] = 16'h2f5b;
mem_array[26236] = 16'h3e03;
mem_array[26239] = 16'h9ed8;
mem_array[26238] = 16'hbf1d;
mem_array[26241] = 16'hc6c3;
mem_array[26240] = 16'h3d54;
mem_array[26243] = 16'hf7d3;
mem_array[26242] = 16'h3d5d;
mem_array[26245] = 16'h5d84;
mem_array[26244] = 16'hbe15;
mem_array[26247] = 16'hc3c7;
mem_array[26246] = 16'h3e2d;
mem_array[26249] = 16'hfe5e;
mem_array[26248] = 16'h3dd2;
mem_array[26251] = 16'he17b;
mem_array[26250] = 16'h3db6;
mem_array[26253] = 16'h07f8;
mem_array[26252] = 16'hbf08;
mem_array[26255] = 16'hde2c;
mem_array[26254] = 16'h3db3;
mem_array[26257] = 16'hfe6a;
mem_array[26256] = 16'h3ecc;
mem_array[26259] = 16'h2b69;
mem_array[26258] = 16'h3e35;
mem_array[26261] = 16'h03bc;
mem_array[26260] = 16'h3e5d;
mem_array[26263] = 16'h09ea;
mem_array[26262] = 16'h3e07;
mem_array[26265] = 16'hc433;
mem_array[26264] = 16'h3e1c;
mem_array[26267] = 16'hc0d2;
mem_array[26266] = 16'hbc97;
mem_array[26269] = 16'ha12b;
mem_array[26268] = 16'h3df5;
mem_array[26271] = 16'h6c65;
mem_array[26270] = 16'h3ef1;
mem_array[26273] = 16'hf6e7;
mem_array[26272] = 16'hbd7e;
mem_array[26275] = 16'h1f52;
mem_array[26274] = 16'h3d1d;
mem_array[26277] = 16'hf8a6;
mem_array[26276] = 16'hbc7c;
mem_array[26279] = 16'hba1a;
mem_array[26278] = 16'h3ec3;
mem_array[26281] = 16'h8a4d;
mem_array[26280] = 16'hbef0;
mem_array[26283] = 16'h956d;
mem_array[26282] = 16'h3e0f;
mem_array[26285] = 16'h824d;
mem_array[26284] = 16'h3dab;
mem_array[26287] = 16'h0e18;
mem_array[26286] = 16'hbd8c;
mem_array[26289] = 16'h7291;
mem_array[26288] = 16'h3e21;
mem_array[26291] = 16'h97f2;
mem_array[26290] = 16'h3e73;
mem_array[26293] = 16'hf29d;
mem_array[26292] = 16'hbe0b;
mem_array[26295] = 16'h0f48;
mem_array[26294] = 16'h3e0f;
mem_array[26297] = 16'h1751;
mem_array[26296] = 16'hbdda;
mem_array[26299] = 16'h731f;
mem_array[26298] = 16'hbf55;
mem_array[26301] = 16'h3e1e;
mem_array[26300] = 16'hbd32;
mem_array[26303] = 16'hf372;
mem_array[26302] = 16'hbd60;
mem_array[26305] = 16'hdd8a;
mem_array[26304] = 16'hbe75;
mem_array[26307] = 16'hba1e;
mem_array[26306] = 16'hbe80;
mem_array[26309] = 16'h4e23;
mem_array[26308] = 16'hbe1d;
mem_array[26311] = 16'h8d0c;
mem_array[26310] = 16'hbd05;
mem_array[26313] = 16'h0d47;
mem_array[26312] = 16'hbfec;
mem_array[26315] = 16'ha7e6;
mem_array[26314] = 16'h3daf;
mem_array[26317] = 16'hdb22;
mem_array[26316] = 16'h3e89;
mem_array[26319] = 16'hb590;
mem_array[26318] = 16'hbc92;
mem_array[26321] = 16'h620b;
mem_array[26320] = 16'h3e77;
mem_array[26323] = 16'h5f20;
mem_array[26322] = 16'h3e22;
mem_array[26325] = 16'h53d4;
mem_array[26324] = 16'hbd63;
mem_array[26327] = 16'h8cb4;
mem_array[26326] = 16'h3dc6;
mem_array[26329] = 16'hab89;
mem_array[26328] = 16'h3e55;
mem_array[26331] = 16'hc9fc;
mem_array[26330] = 16'h3ead;
mem_array[26333] = 16'h8405;
mem_array[26332] = 16'hbecf;
mem_array[26335] = 16'h3b28;
mem_array[26334] = 16'hbcba;
mem_array[26337] = 16'hacf1;
mem_array[26336] = 16'hbe81;
mem_array[26339] = 16'h4468;
mem_array[26338] = 16'hbe67;
mem_array[26341] = 16'h68e4;
mem_array[26340] = 16'hbf1f;
mem_array[26343] = 16'h31a5;
mem_array[26342] = 16'h3e88;
mem_array[26345] = 16'hce74;
mem_array[26344] = 16'h3d83;
mem_array[26347] = 16'h7fdf;
mem_array[26346] = 16'hbe9d;
mem_array[26349] = 16'h28e9;
mem_array[26348] = 16'hbcbd;
mem_array[26351] = 16'h0fa2;
mem_array[26350] = 16'hbc6d;
mem_array[26353] = 16'h527d;
mem_array[26352] = 16'h3d9c;
mem_array[26355] = 16'he798;
mem_array[26354] = 16'h3db6;
mem_array[26357] = 16'hac8b;
mem_array[26356] = 16'h3e75;
mem_array[26359] = 16'hde6a;
mem_array[26358] = 16'hbe49;
mem_array[26361] = 16'haa6f;
mem_array[26360] = 16'hbd95;
mem_array[26363] = 16'hb131;
mem_array[26362] = 16'h3ac1;
mem_array[26365] = 16'h3f63;
mem_array[26364] = 16'h3e9e;
mem_array[26367] = 16'h498d;
mem_array[26366] = 16'h3e47;
mem_array[26369] = 16'h2bda;
mem_array[26368] = 16'h3e04;
mem_array[26371] = 16'h99b0;
mem_array[26370] = 16'h3bfd;
mem_array[26373] = 16'h9774;
mem_array[26372] = 16'hc019;
mem_array[26375] = 16'h6982;
mem_array[26374] = 16'hbca3;
mem_array[26377] = 16'hbc97;
mem_array[26376] = 16'h3e98;
mem_array[26379] = 16'h0e33;
mem_array[26378] = 16'hbb25;
mem_array[26381] = 16'h4f18;
mem_array[26380] = 16'h3e90;
mem_array[26383] = 16'h163b;
mem_array[26382] = 16'h3d0f;
mem_array[26385] = 16'hd884;
mem_array[26384] = 16'h3e8c;
mem_array[26387] = 16'hf34f;
mem_array[26386] = 16'h3e09;
mem_array[26389] = 16'h500f;
mem_array[26388] = 16'h3e8d;
mem_array[26391] = 16'h2299;
mem_array[26390] = 16'h3f15;
mem_array[26393] = 16'he171;
mem_array[26392] = 16'hbdac;
mem_array[26395] = 16'h5884;
mem_array[26394] = 16'hbeec;
mem_array[26397] = 16'hee06;
mem_array[26396] = 16'h3c60;
mem_array[26399] = 16'hfa93;
mem_array[26398] = 16'hbe1e;
mem_array[26401] = 16'h1f96;
mem_array[26400] = 16'hbf40;
mem_array[26403] = 16'h2dd2;
mem_array[26402] = 16'hbd65;
mem_array[26405] = 16'h7277;
mem_array[26404] = 16'hbe8a;
mem_array[26407] = 16'hd983;
mem_array[26406] = 16'hbdf0;
mem_array[26409] = 16'h5f47;
mem_array[26408] = 16'h3d86;
mem_array[26411] = 16'h7f19;
mem_array[26410] = 16'h3c01;
mem_array[26413] = 16'hc1df;
mem_array[26412] = 16'h3ec8;
mem_array[26415] = 16'h9679;
mem_array[26414] = 16'h3ca0;
mem_array[26417] = 16'h3b88;
mem_array[26416] = 16'h3f17;
mem_array[26419] = 16'h7bf6;
mem_array[26418] = 16'hbf1a;
mem_array[26421] = 16'h507e;
mem_array[26420] = 16'h3c96;
mem_array[26423] = 16'h5e54;
mem_array[26422] = 16'hbc11;
mem_array[26425] = 16'h746b;
mem_array[26424] = 16'h3e8a;
mem_array[26427] = 16'hbd85;
mem_array[26426] = 16'hbe1e;
mem_array[26429] = 16'hff17;
mem_array[26428] = 16'h3e25;
mem_array[26431] = 16'he166;
mem_array[26430] = 16'hbbb1;
mem_array[26433] = 16'h1593;
mem_array[26432] = 16'hc012;
mem_array[26435] = 16'h7fc2;
mem_array[26434] = 16'hbe09;
mem_array[26437] = 16'h32fb;
mem_array[26436] = 16'h3f11;
mem_array[26439] = 16'h33c9;
mem_array[26438] = 16'h3e8b;
mem_array[26441] = 16'h9742;
mem_array[26440] = 16'h3dfe;
mem_array[26443] = 16'h9a9d;
mem_array[26442] = 16'h3e50;
mem_array[26445] = 16'h816f;
mem_array[26444] = 16'h3ea2;
mem_array[26447] = 16'h0edf;
mem_array[26446] = 16'h3e4c;
mem_array[26449] = 16'h0b94;
mem_array[26448] = 16'hbcb7;
mem_array[26451] = 16'h3549;
mem_array[26450] = 16'h3dff;
mem_array[26453] = 16'h4b57;
mem_array[26452] = 16'h3e06;
mem_array[26455] = 16'h447a;
mem_array[26454] = 16'hbf71;
mem_array[26457] = 16'hcb0b;
mem_array[26456] = 16'hbd9d;
mem_array[26459] = 16'h861a;
mem_array[26458] = 16'h3e85;
mem_array[26461] = 16'hdc25;
mem_array[26460] = 16'h3e88;
mem_array[26463] = 16'hb726;
mem_array[26462] = 16'h3d86;
mem_array[26465] = 16'hee8e;
mem_array[26464] = 16'hbc47;
mem_array[26467] = 16'ha0d3;
mem_array[26466] = 16'h3e2e;
mem_array[26469] = 16'h56e0;
mem_array[26468] = 16'h3dad;
mem_array[26471] = 16'h13b5;
mem_array[26470] = 16'hbe00;
mem_array[26473] = 16'h66e7;
mem_array[26472] = 16'h3dc9;
mem_array[26475] = 16'h7df0;
mem_array[26474] = 16'hbe06;
mem_array[26477] = 16'hed4b;
mem_array[26476] = 16'h3e13;
mem_array[26479] = 16'haaa7;
mem_array[26478] = 16'hbe4d;
mem_array[26481] = 16'ha98a;
mem_array[26480] = 16'hbd16;
mem_array[26483] = 16'hcc50;
mem_array[26482] = 16'hbd7d;
mem_array[26485] = 16'hc16f;
mem_array[26484] = 16'h3d56;
mem_array[26487] = 16'h4f5e;
mem_array[26486] = 16'h3e77;
mem_array[26489] = 16'h4e8a;
mem_array[26488] = 16'hbd40;
mem_array[26491] = 16'h2348;
mem_array[26490] = 16'hbea4;
mem_array[26493] = 16'h3204;
mem_array[26492] = 16'hbf7f;
mem_array[26495] = 16'h81b6;
mem_array[26494] = 16'h3cb9;
mem_array[26497] = 16'he5b5;
mem_array[26496] = 16'h3ef7;
mem_array[26499] = 16'h36ac;
mem_array[26498] = 16'hbd72;
mem_array[26501] = 16'h41e2;
mem_array[26500] = 16'h3e9a;
mem_array[26503] = 16'h9c54;
mem_array[26502] = 16'h3de9;
mem_array[26505] = 16'hd400;
mem_array[26504] = 16'h3da1;
mem_array[26507] = 16'hb551;
mem_array[26506] = 16'h3b39;
mem_array[26509] = 16'hc16b;
mem_array[26508] = 16'h3f0e;
mem_array[26511] = 16'hfde8;
mem_array[26510] = 16'h3f44;
mem_array[26513] = 16'h1e4a;
mem_array[26512] = 16'h3c89;
mem_array[26515] = 16'h21e3;
mem_array[26514] = 16'hbf84;
mem_array[26517] = 16'hb33b;
mem_array[26516] = 16'hbe4d;
mem_array[26519] = 16'he0a3;
mem_array[26518] = 16'h3e2e;
mem_array[26521] = 16'h057b;
mem_array[26520] = 16'h3ef5;
mem_array[26523] = 16'h4bb7;
mem_array[26522] = 16'h3d91;
mem_array[26525] = 16'h4c65;
mem_array[26524] = 16'hbe40;
mem_array[26527] = 16'hae24;
mem_array[26526] = 16'h3d23;
mem_array[26529] = 16'h6ccc;
mem_array[26528] = 16'h3e7e;
mem_array[26531] = 16'h44e9;
mem_array[26530] = 16'h3e7c;
mem_array[26533] = 16'h06b6;
mem_array[26532] = 16'h3d9f;
mem_array[26535] = 16'h6fa8;
mem_array[26534] = 16'h3dc6;
mem_array[26537] = 16'hd9e8;
mem_array[26536] = 16'h3dbb;
mem_array[26539] = 16'hb566;
mem_array[26538] = 16'hbdef;
mem_array[26541] = 16'hc81f;
mem_array[26540] = 16'hbd91;
mem_array[26543] = 16'h36bb;
mem_array[26542] = 16'hbd9e;
mem_array[26545] = 16'hc874;
mem_array[26544] = 16'h3e59;
mem_array[26547] = 16'h75ca;
mem_array[26546] = 16'hbd5d;
mem_array[26549] = 16'hab4c;
mem_array[26548] = 16'hbcdb;
mem_array[26551] = 16'hd316;
mem_array[26550] = 16'hbd07;
mem_array[26553] = 16'hdad7;
mem_array[26552] = 16'hbf19;
mem_array[26555] = 16'h94e9;
mem_array[26554] = 16'h3dd3;
mem_array[26557] = 16'h589c;
mem_array[26556] = 16'h3ea2;
mem_array[26559] = 16'h9723;
mem_array[26558] = 16'h3db1;
mem_array[26561] = 16'h3376;
mem_array[26560] = 16'h3eaf;
mem_array[26563] = 16'h8e3d;
mem_array[26562] = 16'h3e06;
mem_array[26565] = 16'h8a8e;
mem_array[26564] = 16'h3f47;
mem_array[26567] = 16'h15b2;
mem_array[26566] = 16'h3e82;
mem_array[26569] = 16'hd357;
mem_array[26568] = 16'h3f40;
mem_array[26571] = 16'h5e99;
mem_array[26570] = 16'h3ddf;
mem_array[26573] = 16'h2b79;
mem_array[26572] = 16'hbeb2;
mem_array[26575] = 16'h29bc;
mem_array[26574] = 16'hc007;
mem_array[26577] = 16'h8bf4;
mem_array[26576] = 16'hbe96;
mem_array[26579] = 16'h58ce;
mem_array[26578] = 16'h3ea9;
mem_array[26581] = 16'hcf72;
mem_array[26580] = 16'h3e56;
mem_array[26583] = 16'hcd23;
mem_array[26582] = 16'hbdc9;
mem_array[26585] = 16'hd08b;
mem_array[26584] = 16'hbe9c;
mem_array[26587] = 16'ha60a;
mem_array[26586] = 16'h3e43;
mem_array[26589] = 16'hde28;
mem_array[26588] = 16'h3e89;
mem_array[26591] = 16'h7799;
mem_array[26590] = 16'h3eee;
mem_array[26593] = 16'h9a00;
mem_array[26592] = 16'h3edf;
mem_array[26595] = 16'h8cab;
mem_array[26594] = 16'h3e46;
mem_array[26597] = 16'h8a5f;
mem_array[26596] = 16'h3ed9;
mem_array[26599] = 16'h48e5;
mem_array[26598] = 16'hbdd5;
mem_array[26601] = 16'h6412;
mem_array[26600] = 16'hbde5;
mem_array[26603] = 16'haa5b;
mem_array[26602] = 16'h3dce;
mem_array[26605] = 16'h8f63;
mem_array[26604] = 16'h3db2;
mem_array[26607] = 16'h77ee;
mem_array[26606] = 16'hbea8;
mem_array[26609] = 16'hcc94;
mem_array[26608] = 16'hbe14;
mem_array[26611] = 16'hcb3c;
mem_array[26610] = 16'h3d9f;
mem_array[26613] = 16'ha9c6;
mem_array[26612] = 16'hbde1;
mem_array[26615] = 16'h2411;
mem_array[26614] = 16'hbe7e;
mem_array[26617] = 16'h2394;
mem_array[26616] = 16'hbcca;
mem_array[26619] = 16'h658d;
mem_array[26618] = 16'h3ce6;
mem_array[26621] = 16'hbbb1;
mem_array[26620] = 16'h3e30;
mem_array[26623] = 16'hcd69;
mem_array[26622] = 16'hbd0d;
mem_array[26625] = 16'h9104;
mem_array[26624] = 16'hbe7d;
mem_array[26627] = 16'hc5c2;
mem_array[26626] = 16'h3f06;
mem_array[26629] = 16'h9d75;
mem_array[26628] = 16'h3eee;
mem_array[26631] = 16'h4582;
mem_array[26630] = 16'h3ebf;
mem_array[26633] = 16'hb315;
mem_array[26632] = 16'hbeaf;
mem_array[26635] = 16'h8b74;
mem_array[26634] = 16'hbfd5;
mem_array[26637] = 16'h578d;
mem_array[26636] = 16'hbe03;
mem_array[26639] = 16'h3207;
mem_array[26638] = 16'h3e9d;
mem_array[26641] = 16'he99b;
mem_array[26640] = 16'h3f41;
mem_array[26643] = 16'h318f;
mem_array[26642] = 16'hbf1a;
mem_array[26645] = 16'h4256;
mem_array[26644] = 16'hbada;
mem_array[26647] = 16'h4ee8;
mem_array[26646] = 16'h3f31;
mem_array[26649] = 16'hd4a7;
mem_array[26648] = 16'h3e41;
mem_array[26651] = 16'h5dfc;
mem_array[26650] = 16'hbe28;
mem_array[26653] = 16'h91e6;
mem_array[26652] = 16'h3f47;
mem_array[26655] = 16'h57e9;
mem_array[26654] = 16'h3eb4;
mem_array[26657] = 16'ha24e;
mem_array[26656] = 16'h3ee9;
mem_array[26659] = 16'h9964;
mem_array[26658] = 16'hbc65;
mem_array[26661] = 16'h5d85;
mem_array[26660] = 16'hbdde;
mem_array[26663] = 16'h756f;
mem_array[26662] = 16'h3c08;
mem_array[26665] = 16'h4fc0;
mem_array[26664] = 16'h3e85;
mem_array[26667] = 16'h3e1e;
mem_array[26666] = 16'hbbcd;
mem_array[26669] = 16'h07ff;
mem_array[26668] = 16'h3eee;
mem_array[26671] = 16'h7251;
mem_array[26670] = 16'hbd95;
mem_array[26673] = 16'h1469;
mem_array[26672] = 16'h3f11;
mem_array[26675] = 16'h3af3;
mem_array[26674] = 16'hbe59;
mem_array[26677] = 16'hc129;
mem_array[26676] = 16'hbee2;
mem_array[26679] = 16'h816c;
mem_array[26678] = 16'hbf07;
mem_array[26681] = 16'h9366;
mem_array[26680] = 16'hbf09;
mem_array[26683] = 16'h9151;
mem_array[26682] = 16'h3e16;
mem_array[26685] = 16'h5634;
mem_array[26684] = 16'hbf64;
mem_array[26687] = 16'h5c2b;
mem_array[26686] = 16'h3f10;
mem_array[26689] = 16'h5aa1;
mem_array[26688] = 16'h3f62;
mem_array[26691] = 16'hbfaa;
mem_array[26690] = 16'hbd36;
mem_array[26693] = 16'h25a1;
mem_array[26692] = 16'h3edf;
mem_array[26695] = 16'hb78e;
mem_array[26694] = 16'hbfc2;
mem_array[26697] = 16'hbcfe;
mem_array[26696] = 16'h3ea0;
mem_array[26699] = 16'hf53c;
mem_array[26698] = 16'hbecd;
mem_array[26701] = 16'h052f;
mem_array[26700] = 16'h3eb5;
mem_array[26703] = 16'hcfaa;
mem_array[26702] = 16'h3ec0;
mem_array[26705] = 16'h1c53;
mem_array[26704] = 16'h3e3c;
mem_array[26707] = 16'heb03;
mem_array[26706] = 16'hbd7d;
mem_array[26709] = 16'he737;
mem_array[26708] = 16'h3e9f;
mem_array[26711] = 16'h8088;
mem_array[26710] = 16'hbf29;
mem_array[26713] = 16'h2bc9;
mem_array[26712] = 16'h3fa5;
mem_array[26715] = 16'hc396;
mem_array[26714] = 16'h3e5d;
mem_array[26717] = 16'h0e88;
mem_array[26716] = 16'h3f21;
mem_array[26719] = 16'he74d;
mem_array[26718] = 16'h3ed8;
mem_array[26721] = 16'hedb8;
mem_array[26720] = 16'hbda5;
mem_array[26723] = 16'h334b;
mem_array[26722] = 16'h3dc7;
mem_array[26725] = 16'h8164;
mem_array[26724] = 16'h3eef;
mem_array[26727] = 16'h31b2;
mem_array[26726] = 16'h3e75;
mem_array[26729] = 16'hf5da;
mem_array[26728] = 16'h3e8b;
mem_array[26731] = 16'h3119;
mem_array[26730] = 16'h3e2b;
mem_array[26733] = 16'h5c60;
mem_array[26732] = 16'h3f07;
mem_array[26735] = 16'habc6;
mem_array[26734] = 16'hbd05;
mem_array[26737] = 16'h4aed;
mem_array[26736] = 16'hbf3b;
mem_array[26739] = 16'h521d;
mem_array[26738] = 16'h3e8c;
mem_array[26741] = 16'haf39;
mem_array[26740] = 16'hbe90;
mem_array[26743] = 16'h8494;
mem_array[26742] = 16'hbe34;
mem_array[26745] = 16'he13b;
mem_array[26744] = 16'hbf5a;
mem_array[26747] = 16'h2e90;
mem_array[26746] = 16'h3f71;
mem_array[26749] = 16'h8a19;
mem_array[26748] = 16'h3e12;
mem_array[26751] = 16'hf150;
mem_array[26750] = 16'h3da5;
mem_array[26753] = 16'h6574;
mem_array[26752] = 16'h3e2b;
mem_array[26755] = 16'h510d;
mem_array[26754] = 16'hbeba;
mem_array[26757] = 16'h2de5;
mem_array[26756] = 16'h3f01;
mem_array[26759] = 16'h01ff;
mem_array[26758] = 16'h3ddc;
mem_array[26761] = 16'h4306;
mem_array[26760] = 16'hbf48;
mem_array[26763] = 16'h4e7c;
mem_array[26762] = 16'hbd12;
mem_array[26765] = 16'h1c78;
mem_array[26764] = 16'h3f3b;
mem_array[26767] = 16'h82c8;
mem_array[26766] = 16'hbf86;
mem_array[26769] = 16'h69f6;
mem_array[26768] = 16'h3d6f;
mem_array[26771] = 16'h90dc;
mem_array[26770] = 16'hbeda;
mem_array[26773] = 16'h690a;
mem_array[26772] = 16'h3f7c;
mem_array[26775] = 16'h4650;
mem_array[26774] = 16'h3efe;
mem_array[26777] = 16'h17b5;
mem_array[26776] = 16'h3f6d;
mem_array[26779] = 16'hd62d;
mem_array[26778] = 16'h3f80;
mem_array[26781] = 16'h0aeb;
mem_array[26780] = 16'h3d02;
mem_array[26783] = 16'hf864;
mem_array[26782] = 16'h3d99;
mem_array[26785] = 16'h9b91;
mem_array[26784] = 16'h3e28;
mem_array[26787] = 16'h397e;
mem_array[26786] = 16'h3f3e;
mem_array[26789] = 16'h15fd;
mem_array[26788] = 16'h3e5b;
mem_array[26791] = 16'h26a3;
mem_array[26790] = 16'hbe82;
mem_array[26793] = 16'hcf43;
mem_array[26792] = 16'h3fb4;
mem_array[26795] = 16'h90ed;
mem_array[26794] = 16'hbf21;
mem_array[26797] = 16'hee2f;
mem_array[26796] = 16'hbfa1;
mem_array[26799] = 16'h9f16;
mem_array[26798] = 16'h3d25;
mem_array[26801] = 16'h2667;
mem_array[26800] = 16'hbeea;
mem_array[26803] = 16'h5009;
mem_array[26802] = 16'hbf54;
mem_array[26805] = 16'h8503;
mem_array[26804] = 16'hbf7a;
mem_array[26807] = 16'h0d6d;
mem_array[26806] = 16'h3ebf;
mem_array[26809] = 16'h171a;
mem_array[26808] = 16'h3f37;
mem_array[26811] = 16'h554e;
mem_array[26810] = 16'h3ed6;
mem_array[26813] = 16'h85dc;
mem_array[26812] = 16'hbe9b;
mem_array[26815] = 16'h73e2;
mem_array[26814] = 16'hbdd8;
mem_array[26817] = 16'h4ab3;
mem_array[26816] = 16'h3fa0;
mem_array[26819] = 16'h7be6;
mem_array[26818] = 16'h3e76;
mem_array[26821] = 16'he09d;
mem_array[26820] = 16'hbd62;
mem_array[26823] = 16'h22a2;
mem_array[26822] = 16'h3c8e;
mem_array[26825] = 16'h1765;
mem_array[26824] = 16'h3f69;
mem_array[26827] = 16'h2646;
mem_array[26826] = 16'hbecd;
mem_array[26829] = 16'hdeb2;
mem_array[26828] = 16'hbe0c;
mem_array[26831] = 16'h3249;
mem_array[26830] = 16'hbdc4;
mem_array[26833] = 16'h1ddf;
mem_array[26832] = 16'h3fa2;
mem_array[26835] = 16'h3910;
mem_array[26834] = 16'h3f2e;
mem_array[26837] = 16'h2cce;
mem_array[26836] = 16'h3fab;
mem_array[26839] = 16'hf86d;
mem_array[26838] = 16'h3de8;
mem_array[26841] = 16'h8daf;
mem_array[26840] = 16'h3d36;
mem_array[26843] = 16'h65ab;
mem_array[26842] = 16'hbaf1;
mem_array[26845] = 16'h90ac;
mem_array[26844] = 16'hbea2;
mem_array[26847] = 16'h105f;
mem_array[26846] = 16'h3f38;
mem_array[26849] = 16'h2236;
mem_array[26848] = 16'h3da5;
mem_array[26851] = 16'h09ee;
mem_array[26850] = 16'hbd91;
mem_array[26853] = 16'hbbca;
mem_array[26852] = 16'h3f49;
mem_array[26855] = 16'he4f6;
mem_array[26854] = 16'h3d11;
mem_array[26857] = 16'hffd8;
mem_array[26856] = 16'hbc75;
mem_array[26859] = 16'h67bc;
mem_array[26858] = 16'hbecc;
mem_array[26861] = 16'h4cbe;
mem_array[26860] = 16'hbd84;
mem_array[26863] = 16'h2f93;
mem_array[26862] = 16'hbf04;
mem_array[26865] = 16'h4118;
mem_array[26864] = 16'hbe59;
mem_array[26867] = 16'h1b7d;
mem_array[26866] = 16'hbfa1;
mem_array[26869] = 16'hf57c;
mem_array[26868] = 16'h3ef0;
mem_array[26871] = 16'h63b0;
mem_array[26870] = 16'hbafd;
mem_array[26873] = 16'h809b;
mem_array[26872] = 16'h3f98;
mem_array[26875] = 16'hee07;
mem_array[26874] = 16'hbd76;
mem_array[26877] = 16'hd92a;
mem_array[26876] = 16'h3f30;
mem_array[26879] = 16'hccb1;
mem_array[26878] = 16'hbf4d;
mem_array[26881] = 16'h0081;
mem_array[26880] = 16'hbd13;
mem_array[26883] = 16'h38a2;
mem_array[26882] = 16'h3d05;
mem_array[26885] = 16'hacbf;
mem_array[26884] = 16'hbd98;
mem_array[26887] = 16'h7816;
mem_array[26886] = 16'h3c80;
mem_array[26889] = 16'h19a9;
mem_array[26888] = 16'h3d04;
mem_array[26891] = 16'h92fa;
mem_array[26890] = 16'hbd04;
mem_array[26893] = 16'h82ea;
mem_array[26892] = 16'hbd98;
mem_array[26895] = 16'hef2a;
mem_array[26894] = 16'h3da0;
mem_array[26897] = 16'hb172;
mem_array[26896] = 16'hbd16;
mem_array[26899] = 16'he507;
mem_array[26898] = 16'h3c61;
mem_array[26901] = 16'h41bc;
mem_array[26900] = 16'hbba2;
mem_array[26903] = 16'h5bf7;
mem_array[26902] = 16'hbd18;
mem_array[26905] = 16'h4a65;
mem_array[26904] = 16'h3cf1;
mem_array[26907] = 16'h09e1;
mem_array[26906] = 16'h3c94;
mem_array[26909] = 16'hea7e;
mem_array[26908] = 16'h3db2;
mem_array[26911] = 16'h0ac2;
mem_array[26910] = 16'h3c9e;
mem_array[26913] = 16'h056d;
mem_array[26912] = 16'h3cd7;
mem_array[26915] = 16'hb6d9;
mem_array[26914] = 16'h3d53;
mem_array[26917] = 16'h547d;
mem_array[26916] = 16'hbdb3;
mem_array[26919] = 16'h49b1;
mem_array[26918] = 16'hbcac;
mem_array[26921] = 16'hab99;
mem_array[26920] = 16'hbc94;
mem_array[26923] = 16'h398e;
mem_array[26922] = 16'h3e2f;
mem_array[26925] = 16'h6ac3;
mem_array[26924] = 16'hbc35;
mem_array[26927] = 16'h01b0;
mem_array[26926] = 16'h3ac3;
mem_array[26929] = 16'hb6c9;
mem_array[26928] = 16'h3bcc;
mem_array[26931] = 16'h44ab;
mem_array[26930] = 16'h3cec;
mem_array[26933] = 16'h3ea3;
mem_array[26932] = 16'h3db7;
mem_array[26935] = 16'h86b8;
mem_array[26934] = 16'hbcce;
mem_array[26937] = 16'hb5b6;
mem_array[26936] = 16'h3ddc;
mem_array[26939] = 16'h7c12;
mem_array[26938] = 16'h3dd2;
mem_array[26941] = 16'h7605;
mem_array[26940] = 16'h3d73;
mem_array[26943] = 16'h7550;
mem_array[26942] = 16'hbc2d;
mem_array[26945] = 16'hf13c;
mem_array[26944] = 16'hbd6f;
mem_array[26947] = 16'hdea4;
mem_array[26946] = 16'hbd84;
mem_array[26949] = 16'hbcef;
mem_array[26948] = 16'h3d84;
mem_array[26951] = 16'h33ed;
mem_array[26950] = 16'hbca8;
mem_array[26953] = 16'h44a6;
mem_array[26952] = 16'h3f05;
mem_array[26955] = 16'hc3da;
mem_array[26954] = 16'h3f39;
mem_array[26957] = 16'hf174;
mem_array[26956] = 16'h3dc2;
mem_array[26959] = 16'hcb01;
mem_array[26958] = 16'hbd8f;
mem_array[26961] = 16'hedee;
mem_array[26960] = 16'h3d69;
mem_array[26963] = 16'hc0eb;
mem_array[26962] = 16'hbd5a;
mem_array[26965] = 16'hbc3d;
mem_array[26964] = 16'hbd6f;
mem_array[26967] = 16'h6c60;
mem_array[26966] = 16'hbec2;
mem_array[26969] = 16'h459b;
mem_array[26968] = 16'hbdd0;
mem_array[26971] = 16'h70b4;
mem_array[26970] = 16'hbe2c;
mem_array[26973] = 16'hf163;
mem_array[26972] = 16'hbd4d;
mem_array[26975] = 16'h9ad2;
mem_array[26974] = 16'hbd04;
mem_array[26977] = 16'h118d;
mem_array[26976] = 16'hbd34;
mem_array[26979] = 16'ha120;
mem_array[26978] = 16'hbde4;
mem_array[26981] = 16'ha02f;
mem_array[26980] = 16'hbbfb;
mem_array[26983] = 16'h1d50;
mem_array[26982] = 16'h3e9c;
mem_array[26985] = 16'ha11d;
mem_array[26984] = 16'hbcd7;
mem_array[26987] = 16'hd66f;
mem_array[26986] = 16'hbf6a;
mem_array[26989] = 16'h7007;
mem_array[26988] = 16'h3f76;
mem_array[26991] = 16'hcaf4;
mem_array[26990] = 16'hbd9a;
mem_array[26993] = 16'h7f2b;
mem_array[26992] = 16'h3f0b;
mem_array[26995] = 16'h6c30;
mem_array[26994] = 16'hbc72;
mem_array[26997] = 16'hf610;
mem_array[26996] = 16'h3e98;
mem_array[26999] = 16'h2115;
mem_array[26998] = 16'h3d04;
mem_array[27001] = 16'he751;
mem_array[27000] = 16'h3ec9;
mem_array[27003] = 16'hcc84;
mem_array[27002] = 16'h3e10;
mem_array[27005] = 16'hf199;
mem_array[27004] = 16'h3fb7;
mem_array[27007] = 16'h1309;
mem_array[27006] = 16'hbeb4;
mem_array[27009] = 16'ha935;
mem_array[27008] = 16'hbdc6;
mem_array[27011] = 16'h5502;
mem_array[27010] = 16'h3f11;
mem_array[27013] = 16'hb748;
mem_array[27012] = 16'h3f14;
mem_array[27015] = 16'h5eea;
mem_array[27014] = 16'h3eec;
mem_array[27017] = 16'heba3;
mem_array[27016] = 16'hbce8;
mem_array[27019] = 16'h3504;
mem_array[27018] = 16'hbe28;
mem_array[27021] = 16'hfef0;
mem_array[27020] = 16'hbd4d;
mem_array[27023] = 16'he64c;
mem_array[27022] = 16'h3ca5;
mem_array[27025] = 16'h357c;
mem_array[27024] = 16'hbdea;
mem_array[27027] = 16'h8281;
mem_array[27026] = 16'hbea1;
mem_array[27029] = 16'h5ffa;
mem_array[27028] = 16'h3ec6;
mem_array[27031] = 16'hca27;
mem_array[27030] = 16'hbe8d;
mem_array[27033] = 16'h7380;
mem_array[27032] = 16'h3f1c;
mem_array[27035] = 16'h556a;
mem_array[27034] = 16'hbdf7;
mem_array[27037] = 16'hb958;
mem_array[27036] = 16'hbf8f;
mem_array[27039] = 16'hb170;
mem_array[27038] = 16'h3f2f;
mem_array[27041] = 16'h2efd;
mem_array[27040] = 16'hbe8f;
mem_array[27043] = 16'hf132;
mem_array[27042] = 16'hbeb6;
mem_array[27045] = 16'hf8ee;
mem_array[27044] = 16'hbd8b;
mem_array[27047] = 16'h30f3;
mem_array[27046] = 16'hbf81;
mem_array[27049] = 16'h7efe;
mem_array[27048] = 16'h3f4e;
mem_array[27051] = 16'h32e6;
mem_array[27050] = 16'h3efb;
mem_array[27053] = 16'h4f69;
mem_array[27052] = 16'h3f55;
mem_array[27055] = 16'h8601;
mem_array[27054] = 16'h3e9f;
mem_array[27057] = 16'h37af;
mem_array[27056] = 16'hbef3;
mem_array[27059] = 16'hd509;
mem_array[27058] = 16'h3f64;
mem_array[27061] = 16'h866c;
mem_array[27060] = 16'hbd82;
mem_array[27063] = 16'hee7b;
mem_array[27062] = 16'h3ecb;
mem_array[27065] = 16'h305c;
mem_array[27064] = 16'hbe2d;
mem_array[27067] = 16'ha800;
mem_array[27066] = 16'hbfda;
mem_array[27069] = 16'h08b1;
mem_array[27068] = 16'h3f00;
mem_array[27071] = 16'hcc50;
mem_array[27070] = 16'h3d31;
mem_array[27073] = 16'hbd1d;
mem_array[27072] = 16'hbeb8;
mem_array[27075] = 16'h2aee;
mem_array[27074] = 16'hbe2f;
mem_array[27077] = 16'hb320;
mem_array[27076] = 16'h3ed5;
mem_array[27079] = 16'h8a3a;
mem_array[27078] = 16'h3e4e;
mem_array[27081] = 16'h25bf;
mem_array[27080] = 16'hbdb4;
mem_array[27083] = 16'he331;
mem_array[27082] = 16'h3d5a;
mem_array[27085] = 16'hde68;
mem_array[27084] = 16'h3ce1;
mem_array[27087] = 16'hcf40;
mem_array[27086] = 16'hbd91;
mem_array[27089] = 16'h072e;
mem_array[27088] = 16'hbed6;
mem_array[27091] = 16'h5db8;
mem_array[27090] = 16'h3f53;
mem_array[27093] = 16'h99f4;
mem_array[27092] = 16'hbe74;
mem_array[27095] = 16'h6d4e;
mem_array[27094] = 16'hbea1;
mem_array[27097] = 16'h7da8;
mem_array[27096] = 16'hbf0e;
mem_array[27099] = 16'h9944;
mem_array[27098] = 16'h3da0;
mem_array[27101] = 16'hd298;
mem_array[27100] = 16'hbeea;
mem_array[27103] = 16'h22be;
mem_array[27102] = 16'h3d9b;
mem_array[27105] = 16'h59fc;
mem_array[27104] = 16'hbebe;
mem_array[27107] = 16'h7459;
mem_array[27106] = 16'hbe3f;
mem_array[27109] = 16'h47ba;
mem_array[27108] = 16'h3f5a;
mem_array[27111] = 16'h27cd;
mem_array[27110] = 16'h3f1e;
mem_array[27113] = 16'h2777;
mem_array[27112] = 16'h3f34;
mem_array[27115] = 16'h9f0e;
mem_array[27114] = 16'h3e5b;
mem_array[27117] = 16'he8cf;
mem_array[27116] = 16'hbced;
mem_array[27119] = 16'h556f;
mem_array[27118] = 16'h3e80;
mem_array[27121] = 16'h7342;
mem_array[27120] = 16'hbf42;
mem_array[27123] = 16'hee88;
mem_array[27122] = 16'h3f6a;
mem_array[27125] = 16'hb7c7;
mem_array[27124] = 16'hbf95;
mem_array[27127] = 16'h59e6;
mem_array[27126] = 16'h3f04;
mem_array[27129] = 16'h8127;
mem_array[27128] = 16'h3c64;
mem_array[27131] = 16'ha83a;
mem_array[27130] = 16'hbda8;
mem_array[27133] = 16'he9aa;
mem_array[27132] = 16'hbdaf;
mem_array[27135] = 16'h1b69;
mem_array[27134] = 16'h3ed2;
mem_array[27137] = 16'ha09b;
mem_array[27136] = 16'h3e28;
mem_array[27139] = 16'h4cd2;
mem_array[27138] = 16'hbd8c;
mem_array[27141] = 16'hccff;
mem_array[27140] = 16'hbdad;
mem_array[27143] = 16'h74b4;
mem_array[27142] = 16'h3b8a;
mem_array[27145] = 16'h3895;
mem_array[27144] = 16'h3e2d;
mem_array[27147] = 16'h9494;
mem_array[27146] = 16'h3ebd;
mem_array[27149] = 16'h00b9;
mem_array[27148] = 16'hbf2d;
mem_array[27151] = 16'hc021;
mem_array[27150] = 16'hbd70;
mem_array[27153] = 16'h2a0a;
mem_array[27152] = 16'h3e01;
mem_array[27155] = 16'hf387;
mem_array[27154] = 16'hbeba;
mem_array[27157] = 16'he155;
mem_array[27156] = 16'h3cad;
mem_array[27159] = 16'hc7fb;
mem_array[27158] = 16'hbea7;
mem_array[27161] = 16'h9153;
mem_array[27160] = 16'h3e91;
mem_array[27163] = 16'h66fb;
mem_array[27162] = 16'hbe0d;
mem_array[27165] = 16'h09b4;
mem_array[27164] = 16'hbf07;
mem_array[27167] = 16'h0f51;
mem_array[27166] = 16'h3d1b;
mem_array[27169] = 16'hcb03;
mem_array[27168] = 16'h3f62;
mem_array[27171] = 16'h62e8;
mem_array[27170] = 16'hbdf2;
mem_array[27173] = 16'h2f46;
mem_array[27172] = 16'hbec1;
mem_array[27175] = 16'he68a;
mem_array[27174] = 16'hbcb5;
mem_array[27177] = 16'hcdda;
mem_array[27176] = 16'h3f13;
mem_array[27179] = 16'h5914;
mem_array[27178] = 16'hbe9b;
mem_array[27181] = 16'h669b;
mem_array[27180] = 16'hbf15;
mem_array[27183] = 16'h0806;
mem_array[27182] = 16'h3cd3;
mem_array[27185] = 16'h856b;
mem_array[27184] = 16'hbf8d;
mem_array[27187] = 16'hb7c5;
mem_array[27186] = 16'h3e9f;
mem_array[27189] = 16'h5b5a;
mem_array[27188] = 16'h3e89;
mem_array[27191] = 16'hdd9c;
mem_array[27190] = 16'h3de7;
mem_array[27193] = 16'h9c10;
mem_array[27192] = 16'hbeae;
mem_array[27195] = 16'h6a59;
mem_array[27194] = 16'hbd6d;
mem_array[27197] = 16'h30de;
mem_array[27196] = 16'hbe0a;
mem_array[27199] = 16'h21aa;
mem_array[27198] = 16'hbeb6;
mem_array[27201] = 16'ha094;
mem_array[27200] = 16'hbd6f;
mem_array[27203] = 16'hb080;
mem_array[27202] = 16'h3dde;
mem_array[27205] = 16'hf4a8;
mem_array[27204] = 16'h3dc0;
mem_array[27207] = 16'h865f;
mem_array[27206] = 16'h3e60;
mem_array[27209] = 16'h185e;
mem_array[27208] = 16'hbf26;
mem_array[27211] = 16'h6415;
mem_array[27210] = 16'h3ea3;
mem_array[27213] = 16'hcb7d;
mem_array[27212] = 16'h3e7d;
mem_array[27215] = 16'hc012;
mem_array[27214] = 16'hbe81;
mem_array[27217] = 16'he6a0;
mem_array[27216] = 16'hbdb7;
mem_array[27219] = 16'hdd0d;
mem_array[27218] = 16'hbd90;
mem_array[27221] = 16'h6293;
mem_array[27220] = 16'h3e26;
mem_array[27223] = 16'hc924;
mem_array[27222] = 16'h3dae;
mem_array[27225] = 16'h59e7;
mem_array[27224] = 16'hbf59;
mem_array[27227] = 16'hd337;
mem_array[27226] = 16'h3e54;
mem_array[27229] = 16'hf76a;
mem_array[27228] = 16'h3d37;
mem_array[27231] = 16'h68dd;
mem_array[27230] = 16'hbd9b;
mem_array[27233] = 16'hbb1a;
mem_array[27232] = 16'h3dc8;
mem_array[27235] = 16'hfd76;
mem_array[27234] = 16'h3f07;
mem_array[27237] = 16'h54b7;
mem_array[27236] = 16'h3efb;
mem_array[27239] = 16'h9da3;
mem_array[27238] = 16'h3e85;
mem_array[27241] = 16'h052a;
mem_array[27240] = 16'hbec3;
mem_array[27243] = 16'hf64e;
mem_array[27242] = 16'h3ed0;
mem_array[27245] = 16'hb83d;
mem_array[27244] = 16'hbfca;
mem_array[27247] = 16'h0d4c;
mem_array[27246] = 16'h3eef;
mem_array[27249] = 16'hc4dc;
mem_array[27248] = 16'h3d57;
mem_array[27251] = 16'hd697;
mem_array[27250] = 16'hbf07;
mem_array[27253] = 16'h43a2;
mem_array[27252] = 16'hbef2;
mem_array[27255] = 16'h1aaf;
mem_array[27254] = 16'hbd16;
mem_array[27257] = 16'hb28f;
mem_array[27256] = 16'h3ea9;
mem_array[27259] = 16'heb16;
mem_array[27258] = 16'h3f3d;
mem_array[27261] = 16'h461a;
mem_array[27260] = 16'hbcdd;
mem_array[27263] = 16'he381;
mem_array[27262] = 16'h3d08;
mem_array[27265] = 16'hae72;
mem_array[27264] = 16'h3edf;
mem_array[27267] = 16'h53a3;
mem_array[27266] = 16'h3f0b;
mem_array[27269] = 16'hbadd;
mem_array[27268] = 16'h3e99;
mem_array[27271] = 16'hc8cf;
mem_array[27270] = 16'h3e81;
mem_array[27273] = 16'h2937;
mem_array[27272] = 16'h3f2b;
mem_array[27275] = 16'hbdf8;
mem_array[27274] = 16'h3dbc;
mem_array[27277] = 16'h8294;
mem_array[27276] = 16'h3db0;
mem_array[27279] = 16'h15df;
mem_array[27278] = 16'h3e47;
mem_array[27281] = 16'hfcda;
mem_array[27280] = 16'hbe3a;
mem_array[27283] = 16'h7cb2;
mem_array[27282] = 16'hbdfe;
mem_array[27285] = 16'h0f9a;
mem_array[27284] = 16'h3d9e;
mem_array[27287] = 16'h20d5;
mem_array[27286] = 16'h3e91;
mem_array[27289] = 16'h35c0;
mem_array[27288] = 16'h3e2f;
mem_array[27291] = 16'h1ad3;
mem_array[27290] = 16'hbb20;
mem_array[27293] = 16'ha8c8;
mem_array[27292] = 16'hbd8c;
mem_array[27295] = 16'hd293;
mem_array[27294] = 16'h3e83;
mem_array[27297] = 16'h471b;
mem_array[27296] = 16'h3df7;
mem_array[27299] = 16'h1956;
mem_array[27298] = 16'h3eb9;
mem_array[27301] = 16'h21f4;
mem_array[27300] = 16'hbd24;
mem_array[27303] = 16'h9a3f;
mem_array[27302] = 16'h3eff;
mem_array[27305] = 16'hca7d;
mem_array[27304] = 16'hc00a;
mem_array[27307] = 16'hfe99;
mem_array[27306] = 16'h3f30;
mem_array[27309] = 16'hc527;
mem_array[27308] = 16'h3e1b;
mem_array[27311] = 16'ha1e4;
mem_array[27310] = 16'hbf54;
mem_array[27313] = 16'he7d1;
mem_array[27312] = 16'hbef2;
mem_array[27315] = 16'h3379;
mem_array[27314] = 16'hbee9;
mem_array[27317] = 16'hdea8;
mem_array[27316] = 16'h3e03;
mem_array[27319] = 16'h3365;
mem_array[27318] = 16'h3d90;
mem_array[27321] = 16'hcf72;
mem_array[27320] = 16'hbd45;
mem_array[27323] = 16'hb299;
mem_array[27322] = 16'hbc4e;
mem_array[27325] = 16'hd540;
mem_array[27324] = 16'h3dbf;
mem_array[27327] = 16'h0c25;
mem_array[27326] = 16'h3dfa;
mem_array[27329] = 16'h1201;
mem_array[27328] = 16'h3e1a;
mem_array[27331] = 16'h10d0;
mem_array[27330] = 16'h3e7e;
mem_array[27333] = 16'h9468;
mem_array[27332] = 16'h3f1f;
mem_array[27335] = 16'h0ad3;
mem_array[27334] = 16'h3e60;
mem_array[27337] = 16'hf750;
mem_array[27336] = 16'h3ec5;
mem_array[27339] = 16'h8842;
mem_array[27338] = 16'h3e85;
mem_array[27341] = 16'hfc51;
mem_array[27340] = 16'hbb97;
mem_array[27343] = 16'h06af;
mem_array[27342] = 16'hbd6c;
mem_array[27345] = 16'hb101;
mem_array[27344] = 16'hbb11;
mem_array[27347] = 16'h3681;
mem_array[27346] = 16'h3ecb;
mem_array[27349] = 16'hd31e;
mem_array[27348] = 16'h3e0b;
mem_array[27351] = 16'h29b6;
mem_array[27350] = 16'h3e28;
mem_array[27353] = 16'hc0c5;
mem_array[27352] = 16'hbe0e;
mem_array[27355] = 16'hcfe6;
mem_array[27354] = 16'hbdcb;
mem_array[27357] = 16'ha450;
mem_array[27356] = 16'hb967;
mem_array[27359] = 16'h81ac;
mem_array[27358] = 16'h3f11;
mem_array[27361] = 16'h6e9c;
mem_array[27360] = 16'h3e85;
mem_array[27363] = 16'h8f27;
mem_array[27362] = 16'h3ea3;
mem_array[27365] = 16'h04df;
mem_array[27364] = 16'hbfb2;
mem_array[27367] = 16'h1100;
mem_array[27366] = 16'h3f12;
mem_array[27369] = 16'hdca9;
mem_array[27368] = 16'h3d9b;
mem_array[27371] = 16'h7052;
mem_array[27370] = 16'hbf9c;
mem_array[27373] = 16'h6334;
mem_array[27372] = 16'hbf34;
mem_array[27375] = 16'ha3de;
mem_array[27374] = 16'hbef3;
mem_array[27377] = 16'hc503;
mem_array[27376] = 16'hbe8b;
mem_array[27379] = 16'h93ec;
mem_array[27378] = 16'hbf20;
mem_array[27381] = 16'h4da1;
mem_array[27380] = 16'h3cc0;
mem_array[27383] = 16'he756;
mem_array[27382] = 16'h3d25;
mem_array[27385] = 16'hcf69;
mem_array[27384] = 16'h3e6e;
mem_array[27387] = 16'h18b4;
mem_array[27386] = 16'hbdd3;
mem_array[27389] = 16'he314;
mem_array[27388] = 16'h3eaf;
mem_array[27391] = 16'h7971;
mem_array[27390] = 16'h3e23;
mem_array[27393] = 16'hced2;
mem_array[27392] = 16'h3e4d;
mem_array[27395] = 16'ha6ca;
mem_array[27394] = 16'hbc84;
mem_array[27397] = 16'h72a4;
mem_array[27396] = 16'h3e86;
mem_array[27399] = 16'hf562;
mem_array[27398] = 16'h3ecf;
mem_array[27401] = 16'h597a;
mem_array[27400] = 16'h3e48;
mem_array[27403] = 16'hf951;
mem_array[27402] = 16'h3e0c;
mem_array[27405] = 16'hff00;
mem_array[27404] = 16'h3e46;
mem_array[27407] = 16'h44ab;
mem_array[27406] = 16'h3eb4;
mem_array[27409] = 16'h4cb3;
mem_array[27408] = 16'h3c93;
mem_array[27411] = 16'h8622;
mem_array[27410] = 16'hbe8b;
mem_array[27413] = 16'h8511;
mem_array[27412] = 16'hbde0;
mem_array[27415] = 16'h269a;
mem_array[27414] = 16'h3d06;
mem_array[27417] = 16'h644a;
mem_array[27416] = 16'hbea9;
mem_array[27419] = 16'hf574;
mem_array[27418] = 16'h3ee2;
mem_array[27421] = 16'h59ba;
mem_array[27420] = 16'hbda7;
mem_array[27423] = 16'hadff;
mem_array[27422] = 16'h3e8a;
mem_array[27425] = 16'h3834;
mem_array[27424] = 16'hbdac;
mem_array[27427] = 16'h53d4;
mem_array[27426] = 16'h3f08;
mem_array[27429] = 16'h95d4;
mem_array[27428] = 16'hbe25;
mem_array[27431] = 16'h4975;
mem_array[27430] = 16'hbf3d;
mem_array[27433] = 16'hb610;
mem_array[27432] = 16'hbed7;
mem_array[27435] = 16'h569e;
mem_array[27434] = 16'hbee8;
mem_array[27437] = 16'h8f15;
mem_array[27436] = 16'h3d6f;
mem_array[27439] = 16'h0e5f;
mem_array[27438] = 16'hbd00;
mem_array[27441] = 16'h20e5;
mem_array[27440] = 16'hbcf7;
mem_array[27443] = 16'h6f37;
mem_array[27442] = 16'h3d73;
mem_array[27445] = 16'h1841;
mem_array[27444] = 16'h3e45;
mem_array[27447] = 16'hf132;
mem_array[27446] = 16'h3eca;
mem_array[27449] = 16'h9308;
mem_array[27448] = 16'h3ead;
mem_array[27451] = 16'h000e;
mem_array[27450] = 16'h3da7;
mem_array[27453] = 16'h59ad;
mem_array[27452] = 16'h3e08;
mem_array[27455] = 16'hadbb;
mem_array[27454] = 16'h3e66;
mem_array[27457] = 16'h4fba;
mem_array[27456] = 16'hbd8d;
mem_array[27459] = 16'h782a;
mem_array[27458] = 16'h3eb0;
mem_array[27461] = 16'haf89;
mem_array[27460] = 16'h3db8;
mem_array[27463] = 16'h0679;
mem_array[27462] = 16'hbe39;
mem_array[27465] = 16'ha6b8;
mem_array[27464] = 16'h3e8c;
mem_array[27467] = 16'h314a;
mem_array[27466] = 16'hbd74;
mem_array[27469] = 16'h6406;
mem_array[27468] = 16'h3e65;
mem_array[27471] = 16'h5eac;
mem_array[27470] = 16'hbf44;
mem_array[27473] = 16'haf1e;
mem_array[27472] = 16'h3de3;
mem_array[27475] = 16'h2858;
mem_array[27474] = 16'hbbd3;
mem_array[27477] = 16'h61c1;
mem_array[27476] = 16'hbd7b;
mem_array[27479] = 16'h5dd8;
mem_array[27478] = 16'h3e95;
mem_array[27481] = 16'h0531;
mem_array[27480] = 16'hbebd;
mem_array[27483] = 16'h5930;
mem_array[27482] = 16'h3f4e;
mem_array[27485] = 16'he234;
mem_array[27484] = 16'h3ebd;
mem_array[27487] = 16'h86d4;
mem_array[27486] = 16'h3f0f;
mem_array[27489] = 16'h5962;
mem_array[27488] = 16'hbe0d;
mem_array[27491] = 16'h967d;
mem_array[27490] = 16'hbee1;
mem_array[27493] = 16'h52c9;
mem_array[27492] = 16'hbe55;
mem_array[27495] = 16'hcd07;
mem_array[27494] = 16'hbf42;
mem_array[27497] = 16'h905c;
mem_array[27496] = 16'h3cd0;
mem_array[27499] = 16'hc103;
mem_array[27498] = 16'hbe0d;
mem_array[27501] = 16'h94f9;
mem_array[27500] = 16'hbd82;
mem_array[27503] = 16'h014a;
mem_array[27502] = 16'hbcfe;
mem_array[27505] = 16'hd337;
mem_array[27504] = 16'h3eec;
mem_array[27507] = 16'hb256;
mem_array[27506] = 16'h3dc3;
mem_array[27509] = 16'h7383;
mem_array[27508] = 16'h3ec5;
mem_array[27511] = 16'h320c;
mem_array[27510] = 16'hbba0;
mem_array[27513] = 16'hd2a1;
mem_array[27512] = 16'h3db3;
mem_array[27515] = 16'h4a78;
mem_array[27514] = 16'h3ccf;
mem_array[27517] = 16'ha965;
mem_array[27516] = 16'h3e4b;
mem_array[27519] = 16'h0dd6;
mem_array[27518] = 16'hba84;
mem_array[27521] = 16'hb384;
mem_array[27520] = 16'h3bda;
mem_array[27523] = 16'hb7fd;
mem_array[27522] = 16'h3d91;
mem_array[27525] = 16'h7596;
mem_array[27524] = 16'h3e88;
mem_array[27527] = 16'h29ae;
mem_array[27526] = 16'h3e4f;
mem_array[27529] = 16'h11cc;
mem_array[27528] = 16'h3d84;
mem_array[27531] = 16'he5f9;
mem_array[27530] = 16'hbf0a;
mem_array[27533] = 16'h7608;
mem_array[27532] = 16'h3e13;
mem_array[27535] = 16'h9ca1;
mem_array[27534] = 16'h3e55;
mem_array[27537] = 16'h1bac;
mem_array[27536] = 16'hbe57;
mem_array[27539] = 16'h5a73;
mem_array[27538] = 16'h3e84;
mem_array[27541] = 16'hf8b3;
mem_array[27540] = 16'h3e82;
mem_array[27543] = 16'hb79f;
mem_array[27542] = 16'hbf56;
mem_array[27545] = 16'h5dec;
mem_array[27544] = 16'hbbe0;
mem_array[27547] = 16'h7d8f;
mem_array[27546] = 16'h3ede;
mem_array[27549] = 16'hdeeb;
mem_array[27548] = 16'hbeb1;
mem_array[27551] = 16'h6d64;
mem_array[27550] = 16'hbea5;
mem_array[27553] = 16'h9f61;
mem_array[27552] = 16'hbf76;
mem_array[27555] = 16'h6b4c;
mem_array[27554] = 16'hbf8c;
mem_array[27557] = 16'h6a83;
mem_array[27556] = 16'hbd9c;
mem_array[27559] = 16'hbff7;
mem_array[27558] = 16'h3dae;
mem_array[27561] = 16'h1c4a;
mem_array[27560] = 16'hbd63;
mem_array[27563] = 16'h2a3a;
mem_array[27562] = 16'hbd9d;
mem_array[27565] = 16'h9259;
mem_array[27564] = 16'h3eaa;
mem_array[27567] = 16'hb51d;
mem_array[27566] = 16'h3d94;
mem_array[27569] = 16'hb3c9;
mem_array[27568] = 16'h3eb1;
mem_array[27571] = 16'h5b2e;
mem_array[27570] = 16'h3e24;
mem_array[27573] = 16'he962;
mem_array[27572] = 16'h3e07;
mem_array[27575] = 16'h7bb0;
mem_array[27574] = 16'hbe40;
mem_array[27577] = 16'h78b6;
mem_array[27576] = 16'h3d0b;
mem_array[27579] = 16'h93ab;
mem_array[27578] = 16'hbe93;
mem_array[27581] = 16'h6346;
mem_array[27580] = 16'hbde7;
mem_array[27583] = 16'h4f37;
mem_array[27582] = 16'h3e24;
mem_array[27585] = 16'h890a;
mem_array[27584] = 16'h3db7;
mem_array[27587] = 16'h2c33;
mem_array[27586] = 16'h3e07;
mem_array[27589] = 16'h9f9e;
mem_array[27588] = 16'h3c52;
mem_array[27591] = 16'h8cf5;
mem_array[27590] = 16'hbec1;
mem_array[27593] = 16'h119e;
mem_array[27592] = 16'h3ee5;
mem_array[27595] = 16'h3cdd;
mem_array[27594] = 16'h3e51;
mem_array[27597] = 16'hcaac;
mem_array[27596] = 16'hbecf;
mem_array[27599] = 16'h41db;
mem_array[27598] = 16'h3eae;
mem_array[27601] = 16'h120c;
mem_array[27600] = 16'h3d66;
mem_array[27603] = 16'h30d4;
mem_array[27602] = 16'hc011;
mem_array[27605] = 16'hf265;
mem_array[27604] = 16'hbc64;
mem_array[27607] = 16'h4247;
mem_array[27606] = 16'hbfa2;
mem_array[27609] = 16'h0403;
mem_array[27608] = 16'hbdef;
mem_array[27611] = 16'h3ac3;
mem_array[27610] = 16'hbe07;
mem_array[27613] = 16'hbe21;
mem_array[27612] = 16'hbe55;
mem_array[27615] = 16'h482d;
mem_array[27614] = 16'hbf8f;
mem_array[27617] = 16'hae63;
mem_array[27616] = 16'hbdec;
mem_array[27619] = 16'h5028;
mem_array[27618] = 16'hbe1d;
mem_array[27621] = 16'h1f91;
mem_array[27620] = 16'hbb17;
mem_array[27623] = 16'h8ddf;
mem_array[27622] = 16'hbd1a;
mem_array[27625] = 16'hdd9f;
mem_array[27624] = 16'hbd3e;
mem_array[27627] = 16'hf699;
mem_array[27626] = 16'hbd84;
mem_array[27629] = 16'hfd76;
mem_array[27628] = 16'h3dc9;
mem_array[27631] = 16'hbbdb;
mem_array[27630] = 16'h3e51;
mem_array[27633] = 16'h371c;
mem_array[27632] = 16'h3e42;
mem_array[27635] = 16'h8581;
mem_array[27634] = 16'h3d6f;
mem_array[27637] = 16'h7883;
mem_array[27636] = 16'hbe12;
mem_array[27639] = 16'h19c8;
mem_array[27638] = 16'hbe7f;
mem_array[27641] = 16'hf1a2;
mem_array[27640] = 16'hbaea;
mem_array[27643] = 16'hd5d1;
mem_array[27642] = 16'h3cf6;
mem_array[27645] = 16'h2dc5;
mem_array[27644] = 16'h3e32;
mem_array[27647] = 16'haeb8;
mem_array[27646] = 16'h3e21;
mem_array[27649] = 16'h26b6;
mem_array[27648] = 16'h3f0b;
mem_array[27651] = 16'hdb63;
mem_array[27650] = 16'h3df8;
mem_array[27653] = 16'h01a3;
mem_array[27652] = 16'h3e84;
mem_array[27655] = 16'h2e7b;
mem_array[27654] = 16'h3cd7;
mem_array[27657] = 16'h7143;
mem_array[27656] = 16'hbec6;
mem_array[27659] = 16'hdbbd;
mem_array[27658] = 16'h3ead;
mem_array[27661] = 16'h5617;
mem_array[27660] = 16'h3d2b;
mem_array[27663] = 16'he3ff;
mem_array[27662] = 16'hbf9c;
mem_array[27665] = 16'h9077;
mem_array[27664] = 16'hbe08;
mem_array[27667] = 16'h2c72;
mem_array[27666] = 16'hbf83;
mem_array[27669] = 16'h8bb2;
mem_array[27668] = 16'h3e97;
mem_array[27671] = 16'hdae2;
mem_array[27670] = 16'hbe12;
mem_array[27673] = 16'h5671;
mem_array[27672] = 16'h3e6b;
mem_array[27675] = 16'h599d;
mem_array[27674] = 16'hbf0a;
mem_array[27677] = 16'hbf03;
mem_array[27676] = 16'hbb8d;
mem_array[27679] = 16'had0b;
mem_array[27678] = 16'h3daf;
mem_array[27681] = 16'hfe30;
mem_array[27680] = 16'hbd43;
mem_array[27683] = 16'h9d3d;
mem_array[27682] = 16'h3bed;
mem_array[27685] = 16'hd488;
mem_array[27684] = 16'hbe99;
mem_array[27687] = 16'h6c45;
mem_array[27686] = 16'h3d05;
mem_array[27689] = 16'hc1d9;
mem_array[27688] = 16'h3e6a;
mem_array[27691] = 16'h9749;
mem_array[27690] = 16'h3e64;
mem_array[27693] = 16'h5d4d;
mem_array[27692] = 16'hbdfc;
mem_array[27695] = 16'hd98c;
mem_array[27694] = 16'h3baa;
mem_array[27697] = 16'hd7e8;
mem_array[27696] = 16'hbdf5;
mem_array[27699] = 16'he6a5;
mem_array[27698] = 16'hbd2c;
mem_array[27701] = 16'hce0a;
mem_array[27700] = 16'h3ee1;
mem_array[27703] = 16'h3ca5;
mem_array[27702] = 16'h3e5b;
mem_array[27705] = 16'h20de;
mem_array[27704] = 16'h3e6d;
mem_array[27707] = 16'h9f70;
mem_array[27706] = 16'hbe6a;
mem_array[27709] = 16'he144;
mem_array[27708] = 16'h3e6b;
mem_array[27711] = 16'hb663;
mem_array[27710] = 16'hbe0c;
mem_array[27713] = 16'h528a;
mem_array[27712] = 16'h3e83;
mem_array[27715] = 16'h550c;
mem_array[27714] = 16'hbe44;
mem_array[27717] = 16'hc003;
mem_array[27716] = 16'h3d87;
mem_array[27719] = 16'h4755;
mem_array[27718] = 16'h3e33;
mem_array[27721] = 16'h7737;
mem_array[27720] = 16'hbe06;
mem_array[27723] = 16'hc596;
mem_array[27722] = 16'h3e20;
mem_array[27725] = 16'h6e20;
mem_array[27724] = 16'h3da0;
mem_array[27727] = 16'h1256;
mem_array[27726] = 16'hbfc3;
mem_array[27729] = 16'hff9e;
mem_array[27728] = 16'h3e29;
mem_array[27731] = 16'h3f17;
mem_array[27730] = 16'h3e28;
mem_array[27733] = 16'h888a;
mem_array[27732] = 16'hbe7a;
mem_array[27735] = 16'h7fc5;
mem_array[27734] = 16'hbf19;
mem_array[27737] = 16'hded1;
mem_array[27736] = 16'h3ebe;
mem_array[27739] = 16'hcc15;
mem_array[27738] = 16'h3da6;
mem_array[27741] = 16'h35c7;
mem_array[27740] = 16'hbdb1;
mem_array[27743] = 16'hbb09;
mem_array[27742] = 16'hbac3;
mem_array[27745] = 16'hccc2;
mem_array[27744] = 16'h3de2;
mem_array[27747] = 16'h9773;
mem_array[27746] = 16'h3d7e;
mem_array[27749] = 16'hea44;
mem_array[27748] = 16'h3e42;
mem_array[27751] = 16'h78f4;
mem_array[27750] = 16'h3e59;
mem_array[27753] = 16'hc113;
mem_array[27752] = 16'hbe80;
mem_array[27755] = 16'ha5e2;
mem_array[27754] = 16'hbd55;
mem_array[27757] = 16'hf026;
mem_array[27756] = 16'hbd2e;
mem_array[27759] = 16'h228f;
mem_array[27758] = 16'hbe97;
mem_array[27761] = 16'hba68;
mem_array[27760] = 16'h3e96;
mem_array[27763] = 16'hd7b8;
mem_array[27762] = 16'hbd0c;
mem_array[27765] = 16'hdd57;
mem_array[27764] = 16'hbebe;
mem_array[27767] = 16'hcf78;
mem_array[27766] = 16'hbdc3;
mem_array[27769] = 16'hbc4b;
mem_array[27768] = 16'h3d85;
mem_array[27771] = 16'h844e;
mem_array[27770] = 16'hbda2;
mem_array[27773] = 16'hb10b;
mem_array[27772] = 16'h3e10;
mem_array[27775] = 16'h4d09;
mem_array[27774] = 16'hbe5c;
mem_array[27777] = 16'h277e;
mem_array[27776] = 16'h3e22;
mem_array[27779] = 16'hdf07;
mem_array[27778] = 16'h3cf9;
mem_array[27781] = 16'h233b;
mem_array[27780] = 16'h3da3;
mem_array[27783] = 16'h09f8;
mem_array[27782] = 16'hbdb8;
mem_array[27785] = 16'ha900;
mem_array[27784] = 16'hbe37;
mem_array[27787] = 16'ha6d5;
mem_array[27786] = 16'hbef0;
mem_array[27789] = 16'h4468;
mem_array[27788] = 16'hbe2c;
mem_array[27791] = 16'ha950;
mem_array[27790] = 16'hbe77;
mem_array[27793] = 16'h7962;
mem_array[27792] = 16'hbe73;
mem_array[27795] = 16'ha310;
mem_array[27794] = 16'hbdb6;
mem_array[27797] = 16'hd9e1;
mem_array[27796] = 16'h3eac;
mem_array[27799] = 16'hddbd;
mem_array[27798] = 16'hbc33;
mem_array[27801] = 16'hab8d;
mem_array[27800] = 16'hbbe3;
mem_array[27803] = 16'h9ddb;
mem_array[27802] = 16'hbdab;
mem_array[27805] = 16'h5356;
mem_array[27804] = 16'hbd78;
mem_array[27807] = 16'h7d15;
mem_array[27806] = 16'hbe40;
mem_array[27809] = 16'ha954;
mem_array[27808] = 16'h3c94;
mem_array[27811] = 16'h5651;
mem_array[27810] = 16'h3e6c;
mem_array[27813] = 16'hf427;
mem_array[27812] = 16'hbe10;
mem_array[27815] = 16'h357d;
mem_array[27814] = 16'h3e1f;
mem_array[27817] = 16'h5775;
mem_array[27816] = 16'h3ebe;
mem_array[27819] = 16'h68bd;
mem_array[27818] = 16'hbe89;
mem_array[27821] = 16'hd16c;
mem_array[27820] = 16'h3eb1;
mem_array[27823] = 16'h03a2;
mem_array[27822] = 16'h3ccf;
mem_array[27825] = 16'h705d;
mem_array[27824] = 16'h3e1e;
mem_array[27827] = 16'h83c7;
mem_array[27826] = 16'hbdb5;
mem_array[27829] = 16'h9681;
mem_array[27828] = 16'h3d7d;
mem_array[27831] = 16'h34fd;
mem_array[27830] = 16'hbdab;
mem_array[27833] = 16'h69c0;
mem_array[27832] = 16'hbb63;
mem_array[27835] = 16'h2b3a;
mem_array[27834] = 16'h3deb;
mem_array[27837] = 16'hde48;
mem_array[27836] = 16'h3ecb;
mem_array[27839] = 16'h521a;
mem_array[27838] = 16'h3ead;
mem_array[27841] = 16'h9649;
mem_array[27840] = 16'h3e59;
mem_array[27843] = 16'h9cb9;
mem_array[27842] = 16'hbea8;
mem_array[27845] = 16'h77a5;
mem_array[27844] = 16'h3db0;
mem_array[27847] = 16'h3641;
mem_array[27846] = 16'hbe51;
mem_array[27849] = 16'hee7c;
mem_array[27848] = 16'hbdaa;
mem_array[27851] = 16'h4b95;
mem_array[27850] = 16'hbe07;
mem_array[27853] = 16'h1a8a;
mem_array[27852] = 16'hbdb7;
mem_array[27855] = 16'h3785;
mem_array[27854] = 16'hbe81;
mem_array[27857] = 16'hd703;
mem_array[27856] = 16'h3e93;
mem_array[27859] = 16'h6bd2;
mem_array[27858] = 16'h3e69;
mem_array[27861] = 16'h8fba;
mem_array[27860] = 16'hbd11;
mem_array[27863] = 16'hb64c;
mem_array[27862] = 16'hbd05;
mem_array[27865] = 16'h4214;
mem_array[27864] = 16'h3e35;
mem_array[27867] = 16'hb37f;
mem_array[27866] = 16'h3e09;
mem_array[27869] = 16'h133d;
mem_array[27868] = 16'hbccc;
mem_array[27871] = 16'hdda4;
mem_array[27870] = 16'h3e43;
mem_array[27873] = 16'h6831;
mem_array[27872] = 16'h3e2c;
mem_array[27875] = 16'ha5da;
mem_array[27874] = 16'h3d1d;
mem_array[27877] = 16'h9cc2;
mem_array[27876] = 16'h3e18;
mem_array[27879] = 16'h8693;
mem_array[27878] = 16'h3c32;
mem_array[27881] = 16'h23fd;
mem_array[27880] = 16'h3ea5;
mem_array[27883] = 16'hd03d;
mem_array[27882] = 16'h3d84;
mem_array[27885] = 16'h95fb;
mem_array[27884] = 16'h3dd2;
mem_array[27887] = 16'h3cac;
mem_array[27886] = 16'hbdbc;
mem_array[27889] = 16'h2eee;
mem_array[27888] = 16'hbdca;
mem_array[27891] = 16'h09b2;
mem_array[27890] = 16'h3e1b;
mem_array[27893] = 16'h0e58;
mem_array[27892] = 16'hbe1a;
mem_array[27895] = 16'haacc;
mem_array[27894] = 16'hbd18;
mem_array[27897] = 16'h9c17;
mem_array[27896] = 16'h3e10;
mem_array[27899] = 16'hf9e0;
mem_array[27898] = 16'h3eba;
mem_array[27901] = 16'h67a2;
mem_array[27900] = 16'hbec1;
mem_array[27903] = 16'hf1e5;
mem_array[27902] = 16'h3e85;
mem_array[27905] = 16'hf646;
mem_array[27904] = 16'h3e69;
mem_array[27907] = 16'h7732;
mem_array[27906] = 16'hbe33;
mem_array[27909] = 16'h6d61;
mem_array[27908] = 16'h3e1a;
mem_array[27911] = 16'hbd09;
mem_array[27910] = 16'h3ca5;
mem_array[27913] = 16'hdf7e;
mem_array[27912] = 16'hbd43;
mem_array[27915] = 16'hed90;
mem_array[27914] = 16'h3dd4;
mem_array[27917] = 16'h7a41;
mem_array[27916] = 16'h3ec3;
mem_array[27919] = 16'h3dcb;
mem_array[27918] = 16'hbf28;
mem_array[27921] = 16'hea48;
mem_array[27920] = 16'hbbd4;
mem_array[27923] = 16'h70bc;
mem_array[27922] = 16'h3c06;
mem_array[27925] = 16'h598d;
mem_array[27924] = 16'h3d78;
mem_array[27927] = 16'he19e;
mem_array[27926] = 16'h3de7;
mem_array[27929] = 16'h1228;
mem_array[27928] = 16'hbb2d;
mem_array[27931] = 16'hc2d3;
mem_array[27930] = 16'hbcb5;
mem_array[27933] = 16'ha42c;
mem_array[27932] = 16'hbfca;
mem_array[27935] = 16'h0fc6;
mem_array[27934] = 16'h3d19;
mem_array[27937] = 16'h0f0a;
mem_array[27936] = 16'h3e8b;
mem_array[27939] = 16'h55d4;
mem_array[27938] = 16'h3d98;
mem_array[27941] = 16'h9d8e;
mem_array[27940] = 16'h3ed6;
mem_array[27943] = 16'h1cb1;
mem_array[27942] = 16'h3e72;
mem_array[27945] = 16'h5346;
mem_array[27944] = 16'h3dc3;
mem_array[27947] = 16'hf2ed;
mem_array[27946] = 16'h3d81;
mem_array[27949] = 16'h03fa;
mem_array[27948] = 16'hbc01;
mem_array[27951] = 16'h700d;
mem_array[27950] = 16'h3f02;
mem_array[27953] = 16'hd8d5;
mem_array[27952] = 16'hbea7;
mem_array[27955] = 16'h820f;
mem_array[27954] = 16'hbe60;
mem_array[27957] = 16'ha195;
mem_array[27956] = 16'h3e8a;
mem_array[27959] = 16'h053f;
mem_array[27958] = 16'h3e2c;
mem_array[27961] = 16'h3d42;
mem_array[27960] = 16'hbd15;
mem_array[27963] = 16'h799e;
mem_array[27962] = 16'hbd73;
mem_array[27965] = 16'heffa;
mem_array[27964] = 16'hbd4b;
mem_array[27967] = 16'hcc76;
mem_array[27966] = 16'hbd72;
mem_array[27969] = 16'h7ace;
mem_array[27968] = 16'hbd43;
mem_array[27971] = 16'ha9dc;
mem_array[27970] = 16'hbc51;
mem_array[27973] = 16'hf8d9;
mem_array[27972] = 16'h3e1a;
mem_array[27975] = 16'ha234;
mem_array[27974] = 16'h3de7;
mem_array[27977] = 16'h35f4;
mem_array[27976] = 16'h3e60;
mem_array[27979] = 16'ha2a7;
mem_array[27978] = 16'hbf3d;
mem_array[27981] = 16'hc398;
mem_array[27980] = 16'h3b26;
mem_array[27983] = 16'h2e5d;
mem_array[27982] = 16'hbdb9;
mem_array[27985] = 16'h529a;
mem_array[27984] = 16'hbbb6;
mem_array[27987] = 16'h65ef;
mem_array[27986] = 16'hbe89;
mem_array[27989] = 16'h7f6e;
mem_array[27988] = 16'h3e6e;
mem_array[27991] = 16'heb93;
mem_array[27990] = 16'h3c81;
mem_array[27993] = 16'h8ed2;
mem_array[27992] = 16'hc031;
mem_array[27995] = 16'hb2b9;
mem_array[27994] = 16'hbe27;
mem_array[27997] = 16'ha5b0;
mem_array[27996] = 16'h3dcc;
mem_array[27999] = 16'hc396;
mem_array[27998] = 16'h3c3b;
mem_array[28001] = 16'h0e5d;
mem_array[28000] = 16'h3f06;
mem_array[28003] = 16'hab32;
mem_array[28002] = 16'h3ec5;
mem_array[28005] = 16'hbafb;
mem_array[28004] = 16'h3cfb;
mem_array[28007] = 16'haf37;
mem_array[28006] = 16'h3dc1;
mem_array[28009] = 16'hfd5c;
mem_array[28008] = 16'hbc33;
mem_array[28011] = 16'h595e;
mem_array[28010] = 16'h3de4;
mem_array[28013] = 16'h3dac;
mem_array[28012] = 16'hbe83;
mem_array[28015] = 16'h3931;
mem_array[28014] = 16'hbe2b;
mem_array[28017] = 16'h3a49;
mem_array[28016] = 16'h3dc5;
mem_array[28019] = 16'hf17f;
mem_array[28018] = 16'h3c7c;
mem_array[28021] = 16'hf889;
mem_array[28020] = 16'h3e1c;
mem_array[28023] = 16'he662;
mem_array[28022] = 16'hbd9a;
mem_array[28025] = 16'h01d3;
mem_array[28024] = 16'h3e98;
mem_array[28027] = 16'hb063;
mem_array[28026] = 16'hbe01;
mem_array[28029] = 16'hfe31;
mem_array[28028] = 16'hbc9f;
mem_array[28031] = 16'hd41e;
mem_array[28030] = 16'hbe75;
mem_array[28033] = 16'h832d;
mem_array[28032] = 16'h3e7a;
mem_array[28035] = 16'h65ce;
mem_array[28034] = 16'h3e9b;
mem_array[28037] = 16'hde42;
mem_array[28036] = 16'h3eab;
mem_array[28039] = 16'he42a;
mem_array[28038] = 16'hbd4b;
mem_array[28041] = 16'hefe1;
mem_array[28040] = 16'hbd31;
mem_array[28043] = 16'h59ef;
mem_array[28042] = 16'h3d7e;
mem_array[28045] = 16'h1639;
mem_array[28044] = 16'h3e32;
mem_array[28047] = 16'hebeb;
mem_array[28046] = 16'h3e56;
mem_array[28049] = 16'ha41c;
mem_array[28048] = 16'hbcb9;
mem_array[28051] = 16'h5082;
mem_array[28050] = 16'hbdca;
mem_array[28053] = 16'h8826;
mem_array[28052] = 16'hc016;
mem_array[28055] = 16'h036e;
mem_array[28054] = 16'h3c32;
mem_array[28057] = 16'h4f4f;
mem_array[28056] = 16'h3e2a;
mem_array[28059] = 16'h9bb2;
mem_array[28058] = 16'h3d86;
mem_array[28061] = 16'h176c;
mem_array[28060] = 16'h3e2a;
mem_array[28063] = 16'h0ab2;
mem_array[28062] = 16'h3ec6;
mem_array[28065] = 16'haeab;
mem_array[28064] = 16'hbda8;
mem_array[28067] = 16'h9db9;
mem_array[28066] = 16'hbd76;
mem_array[28069] = 16'h2a04;
mem_array[28068] = 16'h3e89;
mem_array[28071] = 16'h17c5;
mem_array[28070] = 16'h3e2e;
mem_array[28073] = 16'h11c2;
mem_array[28072] = 16'hbd02;
mem_array[28075] = 16'hc20a;
mem_array[28074] = 16'hbb9e;
mem_array[28077] = 16'h2ad5;
mem_array[28076] = 16'h3eb9;
mem_array[28079] = 16'h7c3d;
mem_array[28078] = 16'h3e6f;
mem_array[28081] = 16'h59b4;
mem_array[28080] = 16'hbc9d;
mem_array[28083] = 16'hacee;
mem_array[28082] = 16'hbe9c;
mem_array[28085] = 16'hd345;
mem_array[28084] = 16'hbe54;
mem_array[28087] = 16'hef9f;
mem_array[28086] = 16'h3e42;
mem_array[28089] = 16'hd4d9;
mem_array[28088] = 16'h3e2a;
mem_array[28091] = 16'hb479;
mem_array[28090] = 16'h3e77;
mem_array[28093] = 16'h87b8;
mem_array[28092] = 16'h3ebb;
mem_array[28095] = 16'hf5db;
mem_array[28094] = 16'h3da2;
mem_array[28097] = 16'hcd4b;
mem_array[28096] = 16'h3e9d;
mem_array[28099] = 16'hd53a;
mem_array[28098] = 16'hbe0d;
mem_array[28101] = 16'h3689;
mem_array[28100] = 16'hbd51;
mem_array[28103] = 16'hbd15;
mem_array[28102] = 16'hbd8b;
mem_array[28105] = 16'h0015;
mem_array[28104] = 16'h3eb8;
mem_array[28107] = 16'h68f8;
mem_array[28106] = 16'h3ca3;
mem_array[28109] = 16'h188e;
mem_array[28108] = 16'hbd87;
mem_array[28111] = 16'h1233;
mem_array[28110] = 16'hbe25;
mem_array[28113] = 16'hec02;
mem_array[28112] = 16'hbf8e;
mem_array[28115] = 16'ha872;
mem_array[28114] = 16'hbed2;
mem_array[28117] = 16'h2eaf;
mem_array[28116] = 16'h3e5a;
mem_array[28119] = 16'h99df;
mem_array[28118] = 16'h3e2b;
mem_array[28121] = 16'ha6ec;
mem_array[28120] = 16'h3e65;
mem_array[28123] = 16'ha58d;
mem_array[28122] = 16'h3df2;
mem_array[28125] = 16'h9999;
mem_array[28124] = 16'h3f01;
mem_array[28127] = 16'h46f5;
mem_array[28126] = 16'h3e9e;
mem_array[28129] = 16'h3048;
mem_array[28128] = 16'h3be7;
mem_array[28131] = 16'h5e6c;
mem_array[28130] = 16'hbe34;
mem_array[28133] = 16'h825c;
mem_array[28132] = 16'hbdd8;
mem_array[28135] = 16'h3a46;
mem_array[28134] = 16'hbe7d;
mem_array[28137] = 16'h4f04;
mem_array[28136] = 16'h3e6d;
mem_array[28139] = 16'hb243;
mem_array[28138] = 16'h3f30;
mem_array[28141] = 16'hdc2a;
mem_array[28140] = 16'h3eda;
mem_array[28143] = 16'h8d3a;
mem_array[28142] = 16'hbd0f;
mem_array[28145] = 16'hbf34;
mem_array[28144] = 16'h3e7f;
mem_array[28147] = 16'h21c9;
mem_array[28146] = 16'hbd8e;
mem_array[28149] = 16'h76e3;
mem_array[28148] = 16'hbcb0;
mem_array[28151] = 16'h120e;
mem_array[28150] = 16'h3d9d;
mem_array[28153] = 16'hc6a2;
mem_array[28152] = 16'h3ee9;
mem_array[28155] = 16'had39;
mem_array[28154] = 16'h3dfd;
mem_array[28157] = 16'h081b;
mem_array[28156] = 16'h3e7e;
mem_array[28159] = 16'h224c;
mem_array[28158] = 16'hbe2a;
mem_array[28161] = 16'h7294;
mem_array[28160] = 16'hbcc0;
mem_array[28163] = 16'hc338;
mem_array[28162] = 16'hbce5;
mem_array[28165] = 16'he122;
mem_array[28164] = 16'h3df2;
mem_array[28167] = 16'h038d;
mem_array[28166] = 16'h3e8e;
mem_array[28169] = 16'hd6f8;
mem_array[28168] = 16'h3e3f;
mem_array[28171] = 16'h9c25;
mem_array[28170] = 16'hbdd3;
mem_array[28173] = 16'h1a49;
mem_array[28172] = 16'hbe82;
mem_array[28175] = 16'h9348;
mem_array[28174] = 16'h3abb;
mem_array[28177] = 16'h7a08;
mem_array[28176] = 16'hbe2f;
mem_array[28179] = 16'h4e23;
mem_array[28178] = 16'h3e96;
mem_array[28181] = 16'h38f5;
mem_array[28180] = 16'h3e98;
mem_array[28183] = 16'h1de6;
mem_array[28182] = 16'h3e43;
mem_array[28185] = 16'h7095;
mem_array[28184] = 16'h3e48;
mem_array[28187] = 16'hee27;
mem_array[28186] = 16'hbce6;
mem_array[28189] = 16'hbf57;
mem_array[28188] = 16'h3e81;
mem_array[28191] = 16'h2b00;
mem_array[28190] = 16'h3f30;
mem_array[28193] = 16'hee92;
mem_array[28192] = 16'h3be6;
mem_array[28195] = 16'h3a6f;
mem_array[28194] = 16'hbf82;
mem_array[28197] = 16'h35a8;
mem_array[28196] = 16'h3e56;
mem_array[28199] = 16'h6be5;
mem_array[28198] = 16'h3f2b;
mem_array[28201] = 16'h1b71;
mem_array[28200] = 16'h3ebc;
mem_array[28203] = 16'he337;
mem_array[28202] = 16'hbe88;
mem_array[28205] = 16'h8a84;
mem_array[28204] = 16'hbd3e;
mem_array[28207] = 16'h754d;
mem_array[28206] = 16'h3bd1;
mem_array[28209] = 16'h8432;
mem_array[28208] = 16'h3ebc;
mem_array[28211] = 16'h2c05;
mem_array[28210] = 16'h3e9e;
mem_array[28213] = 16'hc1c0;
mem_array[28212] = 16'h3e6d;
mem_array[28215] = 16'h9922;
mem_array[28214] = 16'h3f42;
mem_array[28217] = 16'h5ae9;
mem_array[28216] = 16'h3e54;
mem_array[28219] = 16'hff6f;
mem_array[28218] = 16'hbd4b;
mem_array[28221] = 16'h8ce1;
mem_array[28220] = 16'hbd5e;
mem_array[28223] = 16'h1f8a;
mem_array[28222] = 16'h3cd2;
mem_array[28225] = 16'h7c74;
mem_array[28224] = 16'h3e17;
mem_array[28227] = 16'hef01;
mem_array[28226] = 16'h3e74;
mem_array[28229] = 16'had7f;
mem_array[28228] = 16'hbd50;
mem_array[28231] = 16'h1034;
mem_array[28230] = 16'hbdab;
mem_array[28233] = 16'h5bb8;
mem_array[28232] = 16'hbe71;
mem_array[28235] = 16'hf6db;
mem_array[28234] = 16'hbe23;
mem_array[28237] = 16'hb79c;
mem_array[28236] = 16'h3d9c;
mem_array[28239] = 16'h8c58;
mem_array[28238] = 16'hbcf9;
mem_array[28241] = 16'h1419;
mem_array[28240] = 16'hbe2a;
mem_array[28243] = 16'h77d5;
mem_array[28242] = 16'h3dea;
mem_array[28245] = 16'hebcd;
mem_array[28244] = 16'h3dcf;
mem_array[28247] = 16'h786f;
mem_array[28246] = 16'hbd9d;
mem_array[28249] = 16'h9197;
mem_array[28248] = 16'hbde5;
mem_array[28251] = 16'h3294;
mem_array[28250] = 16'h3d9a;
mem_array[28253] = 16'h9009;
mem_array[28252] = 16'h3de3;
mem_array[28255] = 16'hcd19;
mem_array[28254] = 16'hbfe4;
mem_array[28257] = 16'h3976;
mem_array[28256] = 16'h3e39;
mem_array[28259] = 16'h10f0;
mem_array[28258] = 16'h3e6e;
mem_array[28261] = 16'h98e0;
mem_array[28260] = 16'hba84;
mem_array[28263] = 16'hde2a;
mem_array[28262] = 16'hbf23;
mem_array[28265] = 16'h75ec;
mem_array[28264] = 16'h3ea6;
mem_array[28267] = 16'h9034;
mem_array[28266] = 16'h3b02;
mem_array[28269] = 16'hf50c;
mem_array[28268] = 16'hbec5;
mem_array[28271] = 16'hb965;
mem_array[28270] = 16'hbe9f;
mem_array[28273] = 16'hc152;
mem_array[28272] = 16'h3f0f;
mem_array[28275] = 16'h69dd;
mem_array[28274] = 16'h3ec6;
mem_array[28277] = 16'h2008;
mem_array[28276] = 16'h3ef0;
mem_array[28279] = 16'h0f37;
mem_array[28278] = 16'h3ea1;
mem_array[28281] = 16'h3f22;
mem_array[28280] = 16'h3d72;
mem_array[28283] = 16'h67bd;
mem_array[28282] = 16'h3de5;
mem_array[28285] = 16'hbba1;
mem_array[28284] = 16'h3d08;
mem_array[28287] = 16'hde5a;
mem_array[28286] = 16'h3e4b;
mem_array[28289] = 16'hfc74;
mem_array[28288] = 16'hbe7d;
mem_array[28291] = 16'h3674;
mem_array[28290] = 16'hbdff;
mem_array[28293] = 16'h9e94;
mem_array[28292] = 16'h3ea4;
mem_array[28295] = 16'h7507;
mem_array[28294] = 16'hbef3;
mem_array[28297] = 16'ha8b9;
mem_array[28296] = 16'h3dbc;
mem_array[28299] = 16'ha077;
mem_array[28298] = 16'hbe38;
mem_array[28301] = 16'he439;
mem_array[28300] = 16'h3ecb;
mem_array[28303] = 16'h7b07;
mem_array[28302] = 16'h3d1b;
mem_array[28305] = 16'h6a57;
mem_array[28304] = 16'hbf0e;
mem_array[28307] = 16'haffa;
mem_array[28306] = 16'h3df2;
mem_array[28309] = 16'h9527;
mem_array[28308] = 16'hbde6;
mem_array[28311] = 16'h374d;
mem_array[28310] = 16'hbe0a;
mem_array[28313] = 16'h0f75;
mem_array[28312] = 16'h3df2;
mem_array[28315] = 16'h5c9b;
mem_array[28314] = 16'hbf7e;
mem_array[28317] = 16'hfc89;
mem_array[28316] = 16'h3dbc;
mem_array[28319] = 16'h73d7;
mem_array[28318] = 16'hbdb4;
mem_array[28321] = 16'h39c1;
mem_array[28320] = 16'h3e52;
mem_array[28323] = 16'h5ae3;
mem_array[28322] = 16'hbf38;
mem_array[28325] = 16'ha156;
mem_array[28324] = 16'h3eeb;
mem_array[28327] = 16'h1b30;
mem_array[28326] = 16'h3d31;
mem_array[28329] = 16'h506c;
mem_array[28328] = 16'hbeba;
mem_array[28331] = 16'h342b;
mem_array[28330] = 16'h3ea4;
mem_array[28333] = 16'h7444;
mem_array[28332] = 16'h3f42;
mem_array[28335] = 16'h2712;
mem_array[28334] = 16'h3ad0;
mem_array[28337] = 16'h8c22;
mem_array[28336] = 16'h3e38;
mem_array[28339] = 16'h96cc;
mem_array[28338] = 16'h3f89;
mem_array[28341] = 16'h5f4e;
mem_array[28340] = 16'h3d83;
mem_array[28343] = 16'h1639;
mem_array[28342] = 16'h3d9a;
mem_array[28345] = 16'h7536;
mem_array[28344] = 16'hbdec;
mem_array[28347] = 16'hc587;
mem_array[28346] = 16'hbe90;
mem_array[28349] = 16'h0ecb;
mem_array[28348] = 16'h3e70;
mem_array[28351] = 16'h9f68;
mem_array[28350] = 16'hbdb5;
mem_array[28353] = 16'h0235;
mem_array[28352] = 16'hbeaf;
mem_array[28355] = 16'hd2db;
mem_array[28354] = 16'h3e8b;
mem_array[28357] = 16'h0e5a;
mem_array[28356] = 16'hbee3;
mem_array[28359] = 16'h00db;
mem_array[28358] = 16'hbde3;
mem_array[28361] = 16'h17b0;
mem_array[28360] = 16'h3eda;
mem_array[28363] = 16'h157f;
mem_array[28362] = 16'h3e02;
mem_array[28365] = 16'hd76f;
mem_array[28364] = 16'h3e65;
mem_array[28367] = 16'h0efc;
mem_array[28366] = 16'h3e2d;
mem_array[28369] = 16'h7de2;
mem_array[28368] = 16'h3e1d;
mem_array[28371] = 16'h9817;
mem_array[28370] = 16'hbf83;
mem_array[28373] = 16'h2817;
mem_array[28372] = 16'h3f18;
mem_array[28375] = 16'h42e8;
mem_array[28374] = 16'hbe9f;
mem_array[28377] = 16'h72e9;
mem_array[28376] = 16'h3dae;
mem_array[28379] = 16'h7a10;
mem_array[28378] = 16'h3e48;
mem_array[28381] = 16'h482c;
mem_array[28380] = 16'hbe91;
mem_array[28383] = 16'h085c;
mem_array[28382] = 16'hbf20;
mem_array[28385] = 16'hbcc8;
mem_array[28384] = 16'h3fa0;
mem_array[28387] = 16'ha8d6;
mem_array[28386] = 16'h3e59;
mem_array[28389] = 16'hc524;
mem_array[28388] = 16'hbef9;
mem_array[28391] = 16'hf720;
mem_array[28390] = 16'hbf97;
mem_array[28393] = 16'hca6b;
mem_array[28392] = 16'h3f97;
mem_array[28395] = 16'h76d0;
mem_array[28394] = 16'h3da7;
mem_array[28397] = 16'hc3e1;
mem_array[28396] = 16'h3f81;
mem_array[28399] = 16'hbedf;
mem_array[28398] = 16'h3f8a;
mem_array[28401] = 16'h0316;
mem_array[28400] = 16'hbb2c;
mem_array[28403] = 16'hd2a4;
mem_array[28402] = 16'hbd73;
mem_array[28405] = 16'hbba9;
mem_array[28404] = 16'h3ee9;
mem_array[28407] = 16'hf8e4;
mem_array[28406] = 16'h3ec0;
mem_array[28409] = 16'h54f3;
mem_array[28408] = 16'h3f40;
mem_array[28411] = 16'hc7a0;
mem_array[28410] = 16'hbec4;
mem_array[28413] = 16'ha598;
mem_array[28412] = 16'h3f38;
mem_array[28415] = 16'h9bed;
mem_array[28414] = 16'h3eb6;
mem_array[28417] = 16'h9273;
mem_array[28416] = 16'hbfed;
mem_array[28419] = 16'h19e8;
mem_array[28418] = 16'h3e08;
mem_array[28421] = 16'hd74a;
mem_array[28420] = 16'hbf17;
mem_array[28423] = 16'hb893;
mem_array[28422] = 16'hbec4;
mem_array[28425] = 16'h6dcf;
mem_array[28424] = 16'hbf65;
mem_array[28427] = 16'h43fd;
mem_array[28426] = 16'h3f40;
mem_array[28429] = 16'hed1e;
mem_array[28428] = 16'h3f93;
mem_array[28431] = 16'hd939;
mem_array[28430] = 16'hbf0b;
mem_array[28433] = 16'h98d3;
mem_array[28432] = 16'hbd21;
mem_array[28435] = 16'hf25c;
mem_array[28434] = 16'hbeaf;
mem_array[28437] = 16'hbb0c;
mem_array[28436] = 16'h3f1c;
mem_array[28439] = 16'h1b19;
mem_array[28438] = 16'h3e3c;
mem_array[28441] = 16'hc7b7;
mem_array[28440] = 16'h3ebd;
mem_array[28443] = 16'hb08a;
mem_array[28442] = 16'hbe04;
mem_array[28445] = 16'h5b10;
mem_array[28444] = 16'h3f8f;
mem_array[28447] = 16'h7fb8;
mem_array[28446] = 16'hbfa7;
mem_array[28449] = 16'h7fa3;
mem_array[28448] = 16'h3f69;
mem_array[28451] = 16'h8abd;
mem_array[28450] = 16'hbe75;
mem_array[28453] = 16'hf42c;
mem_array[28452] = 16'h3f42;
mem_array[28455] = 16'hdb17;
mem_array[28454] = 16'h3e07;
mem_array[28457] = 16'hbdaf;
mem_array[28456] = 16'h3f58;
mem_array[28459] = 16'h8511;
mem_array[28458] = 16'h3f25;
mem_array[28461] = 16'hd3b1;
mem_array[28460] = 16'hbbcd;
mem_array[28463] = 16'h256c;
mem_array[28462] = 16'h3df8;
mem_array[28465] = 16'h5666;
mem_array[28464] = 16'hbd98;
mem_array[28467] = 16'h5aa1;
mem_array[28466] = 16'h3e8e;
mem_array[28469] = 16'h9c4e;
mem_array[28468] = 16'h3e94;
mem_array[28471] = 16'hb41c;
mem_array[28470] = 16'hbe07;
mem_array[28473] = 16'hb689;
mem_array[28472] = 16'h3fc9;
mem_array[28475] = 16'hff8b;
mem_array[28474] = 16'hbe3c;
mem_array[28477] = 16'h8922;
mem_array[28476] = 16'hbf56;
mem_array[28479] = 16'he205;
mem_array[28478] = 16'h3ea5;
mem_array[28481] = 16'h8964;
mem_array[28480] = 16'hbec1;
mem_array[28483] = 16'hffc3;
mem_array[28482] = 16'hbeb3;
mem_array[28485] = 16'he771;
mem_array[28484] = 16'hbf6d;
mem_array[28487] = 16'h836d;
mem_array[28486] = 16'h3ea4;
mem_array[28489] = 16'haa18;
mem_array[28488] = 16'h3e98;
mem_array[28491] = 16'h9027;
mem_array[28490] = 16'h3f33;
mem_array[28493] = 16'h4d89;
mem_array[28492] = 16'h3d8d;
mem_array[28495] = 16'ha795;
mem_array[28494] = 16'hbe92;
mem_array[28497] = 16'hfdb6;
mem_array[28496] = 16'h3f42;
mem_array[28499] = 16'h43f2;
mem_array[28498] = 16'hbe9d;
mem_array[28501] = 16'he245;
mem_array[28500] = 16'hbd07;
mem_array[28503] = 16'h1f27;
mem_array[28502] = 16'h3dc8;
mem_array[28505] = 16'h2ac8;
mem_array[28504] = 16'h3f59;
mem_array[28507] = 16'h277f;
mem_array[28506] = 16'hbf11;
mem_array[28509] = 16'h328d;
mem_array[28508] = 16'hbe37;
mem_array[28511] = 16'hfffc;
mem_array[28510] = 16'hbdc9;
mem_array[28513] = 16'h618a;
mem_array[28512] = 16'h3fc4;
mem_array[28515] = 16'h9d23;
mem_array[28514] = 16'h3f2d;
mem_array[28517] = 16'h2442;
mem_array[28516] = 16'h3fa9;
mem_array[28519] = 16'h297c;
mem_array[28518] = 16'h3e19;
mem_array[28521] = 16'h9205;
mem_array[28520] = 16'hbce3;
mem_array[28523] = 16'h9af6;
mem_array[28522] = 16'hbd84;
mem_array[28525] = 16'h1965;
mem_array[28524] = 16'hbe00;
mem_array[28527] = 16'h89cf;
mem_array[28526] = 16'h3fa0;
mem_array[28529] = 16'hdee6;
mem_array[28528] = 16'h3d66;
mem_array[28531] = 16'h612e;
mem_array[28530] = 16'hbedf;
mem_array[28533] = 16'h292f;
mem_array[28532] = 16'h3f4b;
mem_array[28535] = 16'hf816;
mem_array[28534] = 16'h3d04;
mem_array[28537] = 16'h1220;
mem_array[28536] = 16'hbed8;
mem_array[28539] = 16'h2c35;
mem_array[28538] = 16'hbf08;
mem_array[28541] = 16'h2736;
mem_array[28540] = 16'hbdec;
mem_array[28543] = 16'hb0d8;
mem_array[28542] = 16'hbecf;
mem_array[28545] = 16'hbecd;
mem_array[28544] = 16'hbd74;
mem_array[28547] = 16'h65c0;
mem_array[28546] = 16'hbf70;
mem_array[28549] = 16'h39c0;
mem_array[28548] = 16'h3f82;
mem_array[28551] = 16'h34c7;
mem_array[28550] = 16'hbd27;
mem_array[28553] = 16'hb464;
mem_array[28552] = 16'h3fa1;
mem_array[28555] = 16'headb;
mem_array[28554] = 16'hbe19;
mem_array[28557] = 16'h63f8;
mem_array[28556] = 16'h3f28;
mem_array[28559] = 16'he2ea;
mem_array[28558] = 16'hbf94;
mem_array[28561] = 16'hef55;
mem_array[28560] = 16'h3d64;
mem_array[28563] = 16'h1a87;
mem_array[28562] = 16'hbc86;
mem_array[28565] = 16'h01ee;
mem_array[28564] = 16'h3d96;
mem_array[28567] = 16'h7230;
mem_array[28566] = 16'h3dac;
mem_array[28569] = 16'h51d8;
mem_array[28568] = 16'hbd3c;
mem_array[28571] = 16'ha2cb;
mem_array[28570] = 16'h3d65;
mem_array[28573] = 16'h28f4;
mem_array[28572] = 16'h3d55;
mem_array[28575] = 16'h6d31;
mem_array[28574] = 16'h3dcd;
mem_array[28577] = 16'hc8fb;
mem_array[28576] = 16'hbbef;
mem_array[28579] = 16'hce74;
mem_array[28578] = 16'hbde4;
mem_array[28581] = 16'he3e9;
mem_array[28580] = 16'hbc3b;
mem_array[28583] = 16'h0428;
mem_array[28582] = 16'hbdc2;
mem_array[28585] = 16'hbac5;
mem_array[28584] = 16'hbd8b;
mem_array[28587] = 16'h6e5a;
mem_array[28586] = 16'h3c28;
mem_array[28589] = 16'h8cb1;
mem_array[28588] = 16'h3ca6;
mem_array[28591] = 16'h0157;
mem_array[28590] = 16'h3c7e;
mem_array[28593] = 16'hb61f;
mem_array[28592] = 16'hbba2;
mem_array[28595] = 16'hdac6;
mem_array[28594] = 16'h3ca5;
mem_array[28597] = 16'hee89;
mem_array[28596] = 16'hbc8f;
mem_array[28599] = 16'hf810;
mem_array[28598] = 16'hbcd6;
mem_array[28601] = 16'h064b;
mem_array[28600] = 16'hb9e3;
mem_array[28603] = 16'hfb14;
mem_array[28602] = 16'h3d87;
mem_array[28605] = 16'haa2c;
mem_array[28604] = 16'hbd10;
mem_array[28607] = 16'he90e;
mem_array[28606] = 16'hbd08;
mem_array[28609] = 16'h213a;
mem_array[28608] = 16'hbd5b;
mem_array[28611] = 16'hb8ea;
mem_array[28610] = 16'h3db8;
mem_array[28613] = 16'hc8b0;
mem_array[28612] = 16'hbdca;
mem_array[28615] = 16'h7215;
mem_array[28614] = 16'hbd62;
mem_array[28617] = 16'h5cdc;
mem_array[28616] = 16'h3d93;
mem_array[28619] = 16'h44a2;
mem_array[28618] = 16'h3d7e;
mem_array[28621] = 16'hbc4d;
mem_array[28620] = 16'h3e00;
mem_array[28623] = 16'h2fda;
mem_array[28622] = 16'h3b21;
mem_array[28625] = 16'h6142;
mem_array[28624] = 16'hbdd1;
mem_array[28627] = 16'h4335;
mem_array[28626] = 16'hbd18;
mem_array[28629] = 16'h8648;
mem_array[28628] = 16'hbdbe;
mem_array[28631] = 16'ha41a;
mem_array[28630] = 16'hbd07;
mem_array[28633] = 16'he369;
mem_array[28632] = 16'h3ee5;
mem_array[28635] = 16'h39c0;
mem_array[28634] = 16'h3e8c;
mem_array[28637] = 16'h707d;
mem_array[28636] = 16'h3e1c;
mem_array[28639] = 16'hcd25;
mem_array[28638] = 16'h3b7a;
mem_array[28641] = 16'h42ac;
mem_array[28640] = 16'h3d7c;
mem_array[28643] = 16'h509d;
mem_array[28642] = 16'hbd38;
mem_array[28645] = 16'h9c0d;
mem_array[28644] = 16'hbe9d;
mem_array[28647] = 16'h062a;
mem_array[28646] = 16'hbe64;
mem_array[28649] = 16'hd17d;
mem_array[28648] = 16'hbb48;
mem_array[28651] = 16'h83c2;
mem_array[28650] = 16'hbf0a;
mem_array[28653] = 16'h0693;
mem_array[28652] = 16'h3d44;
mem_array[28655] = 16'h8367;
mem_array[28654] = 16'h3cf1;
mem_array[28657] = 16'he04d;
mem_array[28656] = 16'hbee9;
mem_array[28659] = 16'hdf3b;
mem_array[28658] = 16'h3dee;
mem_array[28661] = 16'h4210;
mem_array[28660] = 16'hbd6f;
mem_array[28663] = 16'h2da0;
mem_array[28662] = 16'h3e7f;
mem_array[28665] = 16'h59b6;
mem_array[28664] = 16'h3c24;
mem_array[28667] = 16'h38fb;
mem_array[28666] = 16'hbf50;
mem_array[28669] = 16'hbfc4;
mem_array[28668] = 16'h3f5f;
mem_array[28671] = 16'h20a8;
mem_array[28670] = 16'hbe1c;
mem_array[28673] = 16'hbece;
mem_array[28672] = 16'h3f22;
mem_array[28675] = 16'h05bb;
mem_array[28674] = 16'hbd36;
mem_array[28677] = 16'h5dde;
mem_array[28676] = 16'h3eb6;
mem_array[28679] = 16'h7f35;
mem_array[28678] = 16'hbca8;
mem_array[28681] = 16'hc0cb;
mem_array[28680] = 16'h3e13;
mem_array[28683] = 16'h51ca;
mem_array[28682] = 16'h3e9f;
mem_array[28685] = 16'h735e;
mem_array[28684] = 16'h3fa4;
mem_array[28687] = 16'h0b24;
mem_array[28686] = 16'hbee1;
mem_array[28689] = 16'h0a9f;
mem_array[28688] = 16'hbe61;
mem_array[28691] = 16'h51ba;
mem_array[28690] = 16'hbe07;
mem_array[28693] = 16'hd2b8;
mem_array[28692] = 16'h3ed8;
mem_array[28695] = 16'h4773;
mem_array[28694] = 16'h3eda;
mem_array[28697] = 16'hc6e5;
mem_array[28696] = 16'hbe3e;
mem_array[28699] = 16'h6d3f;
mem_array[28698] = 16'hbc16;
mem_array[28701] = 16'h261d;
mem_array[28700] = 16'h3ca3;
mem_array[28703] = 16'h42c0;
mem_array[28702] = 16'h3d62;
mem_array[28705] = 16'ha581;
mem_array[28704] = 16'h3e3d;
mem_array[28707] = 16'h6f1f;
mem_array[28706] = 16'hbe0f;
mem_array[28709] = 16'he47b;
mem_array[28708] = 16'h3ec4;
mem_array[28711] = 16'h757b;
mem_array[28710] = 16'hbda8;
mem_array[28713] = 16'h4e3a;
mem_array[28712] = 16'hbebe;
mem_array[28715] = 16'h7842;
mem_array[28714] = 16'hbe14;
mem_array[28717] = 16'h8917;
mem_array[28716] = 16'hbf88;
mem_array[28719] = 16'ha636;
mem_array[28718] = 16'h3f63;
mem_array[28721] = 16'hfee2;
mem_array[28720] = 16'h3cd4;
mem_array[28723] = 16'h63f7;
mem_array[28722] = 16'hbe90;
mem_array[28725] = 16'h385e;
mem_array[28724] = 16'h3dc9;
mem_array[28727] = 16'h5277;
mem_array[28726] = 16'hbf49;
mem_array[28729] = 16'h3182;
mem_array[28728] = 16'h3f61;
mem_array[28731] = 16'h7c40;
mem_array[28730] = 16'h3eb8;
mem_array[28733] = 16'h0f74;
mem_array[28732] = 16'h3dae;
mem_array[28735] = 16'h9feb;
mem_array[28734] = 16'h3eb0;
mem_array[28737] = 16'h2222;
mem_array[28736] = 16'hbf00;
mem_array[28739] = 16'hb94f;
mem_array[28738] = 16'h3f9f;
mem_array[28741] = 16'h0266;
mem_array[28740] = 16'h3f17;
mem_array[28743] = 16'h7cee;
mem_array[28742] = 16'h3eb5;
mem_array[28745] = 16'h57af;
mem_array[28744] = 16'h3ebc;
mem_array[28747] = 16'h6eb3;
mem_array[28746] = 16'hbf89;
mem_array[28749] = 16'h5f14;
mem_array[28748] = 16'h3ead;
mem_array[28751] = 16'he4bb;
mem_array[28750] = 16'hbe32;
mem_array[28753] = 16'heb23;
mem_array[28752] = 16'hbe3e;
mem_array[28755] = 16'hff51;
mem_array[28754] = 16'h3eb4;
mem_array[28757] = 16'h0ffa;
mem_array[28756] = 16'h3f4f;
mem_array[28759] = 16'hdd70;
mem_array[28758] = 16'h3d21;
mem_array[28761] = 16'hc67e;
mem_array[28760] = 16'hbe0c;
mem_array[28763] = 16'he90c;
mem_array[28762] = 16'hbd84;
mem_array[28765] = 16'h25b3;
mem_array[28764] = 16'h3d07;
mem_array[28767] = 16'hf1ed;
mem_array[28766] = 16'h3c02;
mem_array[28769] = 16'ha3ea;
mem_array[28768] = 16'hbb90;
mem_array[28771] = 16'h3d73;
mem_array[28770] = 16'h3f00;
mem_array[28773] = 16'h87f9;
mem_array[28772] = 16'h3e2e;
mem_array[28775] = 16'he51b;
mem_array[28774] = 16'hbeb2;
mem_array[28777] = 16'h192e;
mem_array[28776] = 16'hbfb5;
mem_array[28779] = 16'h94ed;
mem_array[28778] = 16'h3e3e;
mem_array[28781] = 16'h3a40;
mem_array[28780] = 16'hbebf;
mem_array[28783] = 16'h4c22;
mem_array[28782] = 16'h3e78;
mem_array[28785] = 16'h7a9d;
mem_array[28784] = 16'hbe8e;
mem_array[28787] = 16'h6dd9;
mem_array[28786] = 16'hbee3;
mem_array[28789] = 16'hc88f;
mem_array[28788] = 16'h3eed;
mem_array[28791] = 16'h1431;
mem_array[28790] = 16'h3e9f;
mem_array[28793] = 16'he5be;
mem_array[28792] = 16'h3ef1;
mem_array[28795] = 16'hfad2;
mem_array[28794] = 16'h3ed5;
mem_array[28797] = 16'h7c48;
mem_array[28796] = 16'h3dd0;
mem_array[28799] = 16'hd8ae;
mem_array[28798] = 16'hbe8c;
mem_array[28801] = 16'hbe8b;
mem_array[28800] = 16'h3eb1;
mem_array[28803] = 16'h7a0d;
mem_array[28802] = 16'h3e91;
mem_array[28805] = 16'h856e;
mem_array[28804] = 16'hbfa5;
mem_array[28807] = 16'hde07;
mem_array[28806] = 16'h3ecf;
mem_array[28809] = 16'h0fb2;
mem_array[28808] = 16'h3eea;
mem_array[28811] = 16'h9ac1;
mem_array[28810] = 16'h3dcf;
mem_array[28813] = 16'hd3cf;
mem_array[28812] = 16'hbf2d;
mem_array[28815] = 16'he459;
mem_array[28814] = 16'h3e8f;
mem_array[28817] = 16'h42d7;
mem_array[28816] = 16'h3eb3;
mem_array[28819] = 16'h2c5a;
mem_array[28818] = 16'hbc53;
mem_array[28821] = 16'h6887;
mem_array[28820] = 16'hbce3;
mem_array[28823] = 16'h8cb5;
mem_array[28822] = 16'h3cf3;
mem_array[28825] = 16'h9203;
mem_array[28824] = 16'h3cae;
mem_array[28827] = 16'h8781;
mem_array[28826] = 16'h3e63;
mem_array[28829] = 16'h1c01;
mem_array[28828] = 16'h3c8e;
mem_array[28831] = 16'h2694;
mem_array[28830] = 16'hbd09;
mem_array[28833] = 16'h43ec;
mem_array[28832] = 16'h3dbc;
mem_array[28835] = 16'h79fe;
mem_array[28834] = 16'h3e21;
mem_array[28837] = 16'hf710;
mem_array[28836] = 16'hbd0c;
mem_array[28839] = 16'he0ed;
mem_array[28838] = 16'h3e70;
mem_array[28841] = 16'h3ba7;
mem_array[28840] = 16'h3eab;
mem_array[28843] = 16'h73c6;
mem_array[28842] = 16'hbe93;
mem_array[28845] = 16'ha784;
mem_array[28844] = 16'hbf34;
mem_array[28847] = 16'h3c27;
mem_array[28846] = 16'h3d21;
mem_array[28849] = 16'h102b;
mem_array[28848] = 16'h3ce8;
mem_array[28851] = 16'h8d62;
mem_array[28850] = 16'h3e34;
mem_array[28853] = 16'hc154;
mem_array[28852] = 16'hbdb8;
mem_array[28855] = 16'hcab9;
mem_array[28854] = 16'h3e14;
mem_array[28857] = 16'h2540;
mem_array[28856] = 16'h3da7;
mem_array[28859] = 16'h1be5;
mem_array[28858] = 16'hbeed;
mem_array[28861] = 16'h2162;
mem_array[28860] = 16'hbeac;
mem_array[28863] = 16'h5e91;
mem_array[28862] = 16'hbda0;
mem_array[28865] = 16'hd5f8;
mem_array[28864] = 16'hbf80;
mem_array[28867] = 16'ha52f;
mem_array[28866] = 16'h3d84;
mem_array[28869] = 16'h233f;
mem_array[28868] = 16'h3f17;
mem_array[28871] = 16'hb927;
mem_array[28870] = 16'h3e85;
mem_array[28873] = 16'h5a32;
mem_array[28872] = 16'hbe97;
mem_array[28875] = 16'h8af8;
mem_array[28874] = 16'h3e51;
mem_array[28877] = 16'h0dc3;
mem_array[28876] = 16'h3e74;
mem_array[28879] = 16'h198b;
mem_array[28878] = 16'h3f82;
mem_array[28881] = 16'haa65;
mem_array[28880] = 16'h3c83;
mem_array[28883] = 16'he5a1;
mem_array[28882] = 16'h3bfa;
mem_array[28885] = 16'h81ac;
mem_array[28884] = 16'h3c91;
mem_array[28887] = 16'hbea3;
mem_array[28886] = 16'h3dfe;
mem_array[28889] = 16'h4349;
mem_array[28888] = 16'h3dc8;
mem_array[28891] = 16'hc2f2;
mem_array[28890] = 16'h3e97;
mem_array[28893] = 16'ha411;
mem_array[28892] = 16'hbd44;
mem_array[28895] = 16'h58ed;
mem_array[28894] = 16'hbe65;
mem_array[28897] = 16'h737f;
mem_array[28896] = 16'hbd99;
mem_array[28899] = 16'h989b;
mem_array[28898] = 16'hbda8;
mem_array[28901] = 16'h886a;
mem_array[28900] = 16'hbebe;
mem_array[28903] = 16'h94ac;
mem_array[28902] = 16'h3f01;
mem_array[28905] = 16'hf85b;
mem_array[28904] = 16'hbe40;
mem_array[28907] = 16'hf3e2;
mem_array[28906] = 16'h3f1f;
mem_array[28909] = 16'h6d69;
mem_array[28908] = 16'h3dd8;
mem_array[28911] = 16'hfe96;
mem_array[28910] = 16'hbe69;
mem_array[28913] = 16'h0cbb;
mem_array[28912] = 16'h3e26;
mem_array[28915] = 16'hb9f0;
mem_array[28914] = 16'h3f43;
mem_array[28917] = 16'hf8ef;
mem_array[28916] = 16'h3e59;
mem_array[28919] = 16'hfc7b;
mem_array[28918] = 16'hbe7f;
mem_array[28921] = 16'h348b;
mem_array[28920] = 16'hbeac;
mem_array[28923] = 16'h8c54;
mem_array[28922] = 16'hbede;
mem_array[28925] = 16'hb1b8;
mem_array[28924] = 16'hbf8c;
mem_array[28927] = 16'h58c2;
mem_array[28926] = 16'h3e5c;
mem_array[28929] = 16'h6d96;
mem_array[28928] = 16'h3e12;
mem_array[28931] = 16'hfc62;
mem_array[28930] = 16'h3e61;
mem_array[28933] = 16'hedc3;
mem_array[28932] = 16'hbeab;
mem_array[28935] = 16'h3433;
mem_array[28934] = 16'h3e7e;
mem_array[28937] = 16'h9849;
mem_array[28936] = 16'h3f54;
mem_array[28939] = 16'he889;
mem_array[28938] = 16'hbe83;
mem_array[28941] = 16'h0a72;
mem_array[28940] = 16'hbc58;
mem_array[28943] = 16'h1d06;
mem_array[28942] = 16'h3c11;
mem_array[28945] = 16'hf997;
mem_array[28944] = 16'h3e1b;
mem_array[28947] = 16'h9205;
mem_array[28946] = 16'h3f08;
mem_array[28949] = 16'h19dd;
mem_array[28948] = 16'h3eb8;
mem_array[28951] = 16'hfef7;
mem_array[28950] = 16'h3eb3;
mem_array[28953] = 16'hb983;
mem_array[28952] = 16'h3cdd;
mem_array[28955] = 16'h7c23;
mem_array[28954] = 16'hbd85;
mem_array[28957] = 16'hb876;
mem_array[28956] = 16'h3c22;
mem_array[28959] = 16'h6fc7;
mem_array[28958] = 16'h3dd3;
mem_array[28961] = 16'h8b5a;
mem_array[28960] = 16'h3deb;
mem_array[28963] = 16'h98aa;
mem_array[28962] = 16'h3d66;
mem_array[28965] = 16'h65c8;
mem_array[28964] = 16'hbf36;
mem_array[28967] = 16'hbd2e;
mem_array[28966] = 16'h3e10;
mem_array[28969] = 16'h840e;
mem_array[28968] = 16'hbeb8;
mem_array[28971] = 16'hee0e;
mem_array[28970] = 16'hbf88;
mem_array[28973] = 16'h253c;
mem_array[28972] = 16'h3db3;
mem_array[28975] = 16'he23d;
mem_array[28974] = 16'h3e36;
mem_array[28977] = 16'hc257;
mem_array[28976] = 16'h3e9b;
mem_array[28979] = 16'hac3f;
mem_array[28978] = 16'h3e65;
mem_array[28981] = 16'h908a;
mem_array[28980] = 16'hbe32;
mem_array[28983] = 16'h070f;
mem_array[28982] = 16'h3e5f;
mem_array[28985] = 16'he472;
mem_array[28984] = 16'hbf25;
mem_array[28987] = 16'h05e5;
mem_array[28986] = 16'h3ec1;
mem_array[28989] = 16'hf2c1;
mem_array[28988] = 16'hbe43;
mem_array[28991] = 16'h53f0;
mem_array[28990] = 16'hbdbe;
mem_array[28993] = 16'hd79f;
mem_array[28992] = 16'hbe6a;
mem_array[28995] = 16'h7d2b;
mem_array[28994] = 16'h3e34;
mem_array[28997] = 16'h4cc1;
mem_array[28996] = 16'hbe43;
mem_array[28999] = 16'h7119;
mem_array[28998] = 16'h3d3c;
mem_array[29001] = 16'h3884;
mem_array[29000] = 16'h3d32;
mem_array[29003] = 16'h6f5f;
mem_array[29002] = 16'hbdb6;
mem_array[29005] = 16'hd9ef;
mem_array[29004] = 16'h3db4;
mem_array[29007] = 16'hebd1;
mem_array[29006] = 16'hbe2c;
mem_array[29009] = 16'h3973;
mem_array[29008] = 16'hbd3f;
mem_array[29011] = 16'hcb9d;
mem_array[29010] = 16'h3e62;
mem_array[29013] = 16'h2f7b;
mem_array[29012] = 16'hbea2;
mem_array[29015] = 16'hbdfb;
mem_array[29014] = 16'h3e54;
mem_array[29017] = 16'h098f;
mem_array[29016] = 16'h3ee1;
mem_array[29019] = 16'h4664;
mem_array[29018] = 16'h3eb2;
mem_array[29021] = 16'h07a6;
mem_array[29020] = 16'hbea4;
mem_array[29023] = 16'hedbd;
mem_array[29022] = 16'h3e45;
mem_array[29025] = 16'h200a;
mem_array[29024] = 16'h3d57;
mem_array[29027] = 16'h79d6;
mem_array[29026] = 16'h3e96;
mem_array[29029] = 16'h00d3;
mem_array[29028] = 16'hbe8e;
mem_array[29031] = 16'h2a63;
mem_array[29030] = 16'hbf78;
mem_array[29033] = 16'he38c;
mem_array[29032] = 16'h3bd9;
mem_array[29035] = 16'he234;
mem_array[29034] = 16'hbead;
mem_array[29037] = 16'h3ec1;
mem_array[29036] = 16'hbd6e;
mem_array[29039] = 16'h994b;
mem_array[29038] = 16'h3ee2;
mem_array[29041] = 16'hc645;
mem_array[29040] = 16'hbecb;
mem_array[29043] = 16'he9c6;
mem_array[29042] = 16'hbe8a;
mem_array[29045] = 16'h51ae;
mem_array[29044] = 16'hbbc1;
mem_array[29047] = 16'h3c64;
mem_array[29046] = 16'h3f08;
mem_array[29049] = 16'h7410;
mem_array[29048] = 16'hbe66;
mem_array[29051] = 16'hb966;
mem_array[29050] = 16'hbf35;
mem_array[29053] = 16'h2b9a;
mem_array[29052] = 16'h3dd3;
mem_array[29055] = 16'h16af;
mem_array[29054] = 16'h3dc4;
mem_array[29057] = 16'he284;
mem_array[29056] = 16'hbee3;
mem_array[29059] = 16'h782f;
mem_array[29058] = 16'hbdb7;
mem_array[29061] = 16'h4139;
mem_array[29060] = 16'hbd72;
mem_array[29063] = 16'hcf30;
mem_array[29062] = 16'hbc8e;
mem_array[29065] = 16'h165f;
mem_array[29064] = 16'h3d03;
mem_array[29067] = 16'ha3d6;
mem_array[29066] = 16'h3e10;
mem_array[29069] = 16'h3b85;
mem_array[29068] = 16'h3ec0;
mem_array[29071] = 16'h1c57;
mem_array[29070] = 16'h3ed6;
mem_array[29073] = 16'h931a;
mem_array[29072] = 16'hbdb2;
mem_array[29075] = 16'h4653;
mem_array[29074] = 16'hbd84;
mem_array[29077] = 16'hc355;
mem_array[29076] = 16'h3ed8;
mem_array[29079] = 16'h1c09;
mem_array[29078] = 16'h3e8a;
mem_array[29081] = 16'h569e;
mem_array[29080] = 16'h3eb5;
mem_array[29083] = 16'hd29b;
mem_array[29082] = 16'h3d14;
mem_array[29085] = 16'hfd6a;
mem_array[29084] = 16'hbc8b;
mem_array[29087] = 16'h3857;
mem_array[29086] = 16'h3ecf;
mem_array[29089] = 16'hf721;
mem_array[29088] = 16'hbed9;
mem_array[29091] = 16'h825c;
mem_array[29090] = 16'hbfb1;
mem_array[29093] = 16'h31ec;
mem_array[29092] = 16'h3c92;
mem_array[29095] = 16'hf729;
mem_array[29094] = 16'hbf10;
mem_array[29097] = 16'h12cc;
mem_array[29096] = 16'h3d92;
mem_array[29099] = 16'h0d77;
mem_array[29098] = 16'h3e83;
mem_array[29101] = 16'h14c3;
mem_array[29100] = 16'hbe1b;
mem_array[29103] = 16'h5987;
mem_array[29102] = 16'hbe9b;
mem_array[29105] = 16'h9547;
mem_array[29104] = 16'h3f08;
mem_array[29107] = 16'h6048;
mem_array[29106] = 16'h3f1d;
mem_array[29109] = 16'hc723;
mem_array[29108] = 16'hbeb3;
mem_array[29111] = 16'hd9fb;
mem_array[29110] = 16'hbf74;
mem_array[29113] = 16'hbce5;
mem_array[29112] = 16'hbf1e;
mem_array[29115] = 16'hcb34;
mem_array[29114] = 16'hbd2d;
mem_array[29117] = 16'h33ef;
mem_array[29116] = 16'h3e10;
mem_array[29119] = 16'h7652;
mem_array[29118] = 16'h3e6c;
mem_array[29121] = 16'h3971;
mem_array[29120] = 16'hbdc2;
mem_array[29123] = 16'hf97d;
mem_array[29122] = 16'hbcdb;
mem_array[29125] = 16'h102f;
mem_array[29124] = 16'h3e0e;
mem_array[29127] = 16'h1739;
mem_array[29126] = 16'h3e10;
mem_array[29129] = 16'he5f4;
mem_array[29128] = 16'h3e34;
mem_array[29131] = 16'hf482;
mem_array[29130] = 16'h3e93;
mem_array[29133] = 16'hed4c;
mem_array[29132] = 16'hbc35;
mem_array[29135] = 16'h4e55;
mem_array[29134] = 16'hbe44;
mem_array[29137] = 16'h207e;
mem_array[29136] = 16'h3c6b;
mem_array[29139] = 16'h87c3;
mem_array[29138] = 16'h3e23;
mem_array[29141] = 16'hc8ab;
mem_array[29140] = 16'hbd8d;
mem_array[29143] = 16'hdb81;
mem_array[29142] = 16'h3ced;
mem_array[29145] = 16'hfd10;
mem_array[29144] = 16'h3dbd;
mem_array[29147] = 16'h8057;
mem_array[29146] = 16'h3e9a;
mem_array[29149] = 16'he818;
mem_array[29148] = 16'hbe08;
mem_array[29151] = 16'hc2c3;
mem_array[29150] = 16'hbf27;
mem_array[29153] = 16'hb3f6;
mem_array[29152] = 16'h3d8d;
mem_array[29155] = 16'hffef;
mem_array[29154] = 16'hbe49;
mem_array[29157] = 16'h3f1e;
mem_array[29156] = 16'h3e52;
mem_array[29159] = 16'h592c;
mem_array[29158] = 16'h3e74;
mem_array[29161] = 16'hca99;
mem_array[29160] = 16'h3d15;
mem_array[29163] = 16'hcc14;
mem_array[29162] = 16'hbdf9;
mem_array[29165] = 16'h29cb;
mem_array[29164] = 16'h3eb0;
mem_array[29167] = 16'h5ba6;
mem_array[29166] = 16'h3f27;
mem_array[29169] = 16'h7cc0;
mem_array[29168] = 16'h3e5d;
mem_array[29171] = 16'h6ae0;
mem_array[29170] = 16'hbf69;
mem_array[29173] = 16'h01cc;
mem_array[29172] = 16'hbf88;
mem_array[29175] = 16'h6edb;
mem_array[29174] = 16'hbd41;
mem_array[29177] = 16'hd806;
mem_array[29176] = 16'h3e4e;
mem_array[29179] = 16'h12cc;
mem_array[29178] = 16'hbeaa;
mem_array[29181] = 16'hcedd;
mem_array[29180] = 16'hbdc1;
mem_array[29183] = 16'hb56f;
mem_array[29182] = 16'hbda8;
mem_array[29185] = 16'hfbf4;
mem_array[29184] = 16'h3e41;
mem_array[29187] = 16'h6669;
mem_array[29186] = 16'h3e97;
mem_array[29189] = 16'h7fb0;
mem_array[29188] = 16'h3d88;
mem_array[29191] = 16'h22b5;
mem_array[29190] = 16'h3eb4;
mem_array[29193] = 16'hb57f;
mem_array[29192] = 16'hbd6a;
mem_array[29195] = 16'h674f;
mem_array[29194] = 16'hbd93;
mem_array[29197] = 16'ha411;
mem_array[29196] = 16'h3e90;
mem_array[29199] = 16'ha89b;
mem_array[29198] = 16'h3da3;
mem_array[29201] = 16'h82c1;
mem_array[29200] = 16'h3d6a;
mem_array[29203] = 16'he230;
mem_array[29202] = 16'h3c5e;
mem_array[29205] = 16'h0442;
mem_array[29204] = 16'h3eeb;
mem_array[29207] = 16'he6d6;
mem_array[29206] = 16'h3e25;
mem_array[29209] = 16'hf21d;
mem_array[29208] = 16'hbe30;
mem_array[29211] = 16'he60c;
mem_array[29210] = 16'h3ef9;
mem_array[29213] = 16'hf79a;
mem_array[29212] = 16'hbd5b;
mem_array[29215] = 16'h0fae;
mem_array[29214] = 16'h3e1b;
mem_array[29217] = 16'h9163;
mem_array[29216] = 16'h3e24;
mem_array[29219] = 16'he52b;
mem_array[29218] = 16'h3f0f;
mem_array[29221] = 16'h4b11;
mem_array[29220] = 16'h3e80;
mem_array[29223] = 16'h68c9;
mem_array[29222] = 16'hbfb0;
mem_array[29225] = 16'ha80d;
mem_array[29224] = 16'h3e85;
mem_array[29227] = 16'h5f33;
mem_array[29226] = 16'hbe6c;
mem_array[29229] = 16'h5b53;
mem_array[29228] = 16'hbda9;
mem_array[29231] = 16'hef41;
mem_array[29230] = 16'hbf6e;
mem_array[29233] = 16'h2ff4;
mem_array[29232] = 16'hbfbf;
mem_array[29235] = 16'h7243;
mem_array[29234] = 16'hbea3;
mem_array[29237] = 16'h4161;
mem_array[29236] = 16'h3e09;
mem_array[29239] = 16'hfd2d;
mem_array[29238] = 16'hbe92;
mem_array[29241] = 16'h79e7;
mem_array[29240] = 16'hbd92;
mem_array[29243] = 16'h126b;
mem_array[29242] = 16'h3c49;
mem_array[29245] = 16'hbb8f;
mem_array[29244] = 16'h3e97;
mem_array[29247] = 16'h7abc;
mem_array[29246] = 16'h3dec;
mem_array[29249] = 16'h30e8;
mem_array[29248] = 16'h3e05;
mem_array[29251] = 16'h2ed3;
mem_array[29250] = 16'h3c4a;
mem_array[29253] = 16'h8a4a;
mem_array[29252] = 16'h3d1f;
mem_array[29255] = 16'h5f54;
mem_array[29254] = 16'h3bdc;
mem_array[29257] = 16'hcf09;
mem_array[29256] = 16'hbc99;
mem_array[29259] = 16'h25d3;
mem_array[29258] = 16'hbe90;
mem_array[29261] = 16'h4c19;
mem_array[29260] = 16'hbeb6;
mem_array[29263] = 16'h6784;
mem_array[29262] = 16'h3c85;
mem_array[29265] = 16'heb6c;
mem_array[29264] = 16'h3e16;
mem_array[29267] = 16'h771d;
mem_array[29266] = 16'h3dfd;
mem_array[29269] = 16'h1ef8;
mem_array[29268] = 16'hbde0;
mem_array[29271] = 16'h3772;
mem_array[29270] = 16'h3e1d;
mem_array[29273] = 16'h9b4f;
mem_array[29272] = 16'h3e6d;
mem_array[29275] = 16'h4205;
mem_array[29274] = 16'h3e72;
mem_array[29277] = 16'h8f1a;
mem_array[29276] = 16'h3dbb;
mem_array[29279] = 16'h51a4;
mem_array[29278] = 16'h3df8;
mem_array[29281] = 16'hfec0;
mem_array[29280] = 16'h3ed6;
mem_array[29283] = 16'h5634;
mem_array[29282] = 16'hbff2;
mem_array[29285] = 16'hc6d6;
mem_array[29284] = 16'h3d9d;
mem_array[29287] = 16'h6495;
mem_array[29286] = 16'hbf8a;
mem_array[29289] = 16'h88a5;
mem_array[29288] = 16'h3de4;
mem_array[29291] = 16'h1018;
mem_array[29290] = 16'hbece;
mem_array[29293] = 16'h71eb;
mem_array[29292] = 16'hbfc7;
mem_array[29295] = 16'h4107;
mem_array[29294] = 16'hbef0;
mem_array[29297] = 16'hee40;
mem_array[29296] = 16'h3d5e;
mem_array[29299] = 16'h7c19;
mem_array[29298] = 16'hbda8;
mem_array[29301] = 16'h0712;
mem_array[29300] = 16'hbc33;
mem_array[29303] = 16'hacb0;
mem_array[29302] = 16'hbd0b;
mem_array[29305] = 16'h37ba;
mem_array[29304] = 16'h3e1c;
mem_array[29307] = 16'h1efd;
mem_array[29306] = 16'h3e51;
mem_array[29309] = 16'hec4f;
mem_array[29308] = 16'h3dcc;
mem_array[29311] = 16'h4c70;
mem_array[29310] = 16'h3e1e;
mem_array[29313] = 16'hac71;
mem_array[29312] = 16'h3df3;
mem_array[29315] = 16'h7c44;
mem_array[29314] = 16'h3d07;
mem_array[29317] = 16'hdbca;
mem_array[29316] = 16'hbe75;
mem_array[29319] = 16'hacd9;
mem_array[29318] = 16'h3d1a;
mem_array[29321] = 16'h7742;
mem_array[29320] = 16'hbe82;
mem_array[29323] = 16'hfcbb;
mem_array[29322] = 16'h3d7a;
mem_array[29325] = 16'h1c2a;
mem_array[29324] = 16'h3ed8;
mem_array[29327] = 16'h1a65;
mem_array[29326] = 16'h3e8e;
mem_array[29329] = 16'hc41c;
mem_array[29328] = 16'h3e3d;
mem_array[29331] = 16'h0d26;
mem_array[29330] = 16'hbe9c;
mem_array[29333] = 16'he969;
mem_array[29332] = 16'h3f05;
mem_array[29335] = 16'hb2c8;
mem_array[29334] = 16'h3dda;
mem_array[29337] = 16'h5503;
mem_array[29336] = 16'h3d2f;
mem_array[29339] = 16'h7c60;
mem_array[29338] = 16'hbef2;
mem_array[29341] = 16'h5b72;
mem_array[29340] = 16'h3e13;
mem_array[29343] = 16'h6d17;
mem_array[29342] = 16'hbef7;
mem_array[29345] = 16'h1636;
mem_array[29344] = 16'h3e23;
mem_array[29347] = 16'hbb7f;
mem_array[29346] = 16'hbf5f;
mem_array[29349] = 16'h286c;
mem_array[29348] = 16'h3e93;
mem_array[29351] = 16'h1f71;
mem_array[29350] = 16'hbebb;
mem_array[29353] = 16'h68c1;
mem_array[29352] = 16'hbf6e;
mem_array[29355] = 16'hc171;
mem_array[29354] = 16'hbeef;
mem_array[29357] = 16'hd47c;
mem_array[29356] = 16'h3e02;
mem_array[29359] = 16'h4e41;
mem_array[29358] = 16'h3eb2;
mem_array[29361] = 16'h67af;
mem_array[29360] = 16'hbd9e;
mem_array[29363] = 16'h9c1b;
mem_array[29362] = 16'h3c90;
mem_array[29365] = 16'h99f8;
mem_array[29364] = 16'hbc88;
mem_array[29367] = 16'h189f;
mem_array[29366] = 16'h3ea6;
mem_array[29369] = 16'haeb1;
mem_array[29368] = 16'hbe23;
mem_array[29371] = 16'h37d4;
mem_array[29370] = 16'h3ee4;
mem_array[29373] = 16'ha70c;
mem_array[29372] = 16'hbd3d;
mem_array[29375] = 16'h57e5;
mem_array[29374] = 16'h3e2d;
mem_array[29377] = 16'h30ea;
mem_array[29376] = 16'hbe62;
mem_array[29379] = 16'h6369;
mem_array[29378] = 16'h3e11;
mem_array[29381] = 16'h001b;
mem_array[29380] = 16'h3e0a;
mem_array[29383] = 16'h5b9a;
mem_array[29382] = 16'h3e8d;
mem_array[29385] = 16'ha271;
mem_array[29384] = 16'h3dd3;
mem_array[29387] = 16'h8f3b;
mem_array[29386] = 16'hbe59;
mem_array[29389] = 16'h2b6f;
mem_array[29388] = 16'h3ea1;
mem_array[29391] = 16'h5531;
mem_array[29390] = 16'h3e04;
mem_array[29393] = 16'hb9bf;
mem_array[29392] = 16'h3e9b;
mem_array[29395] = 16'h6885;
mem_array[29394] = 16'hbe30;
mem_array[29397] = 16'h40e4;
mem_array[29396] = 16'h3e7d;
mem_array[29399] = 16'hd35b;
mem_array[29398] = 16'h3e65;
mem_array[29401] = 16'h4a06;
mem_array[29400] = 16'h3d8a;
mem_array[29403] = 16'h7ba2;
mem_array[29402] = 16'h3e9f;
mem_array[29405] = 16'h606f;
mem_array[29404] = 16'h3eac;
mem_array[29407] = 16'hf3fd;
mem_array[29406] = 16'hbf5f;
mem_array[29409] = 16'heaf7;
mem_array[29408] = 16'h3c06;
mem_array[29411] = 16'h74c7;
mem_array[29410] = 16'h3d1b;
mem_array[29413] = 16'h7783;
mem_array[29412] = 16'hbf57;
mem_array[29415] = 16'h3393;
mem_array[29414] = 16'hbeed;
mem_array[29417] = 16'h8ab9;
mem_array[29416] = 16'h3d89;
mem_array[29419] = 16'h039b;
mem_array[29418] = 16'h3f01;
mem_array[29421] = 16'he9d1;
mem_array[29420] = 16'h3ca8;
mem_array[29423] = 16'h9d33;
mem_array[29422] = 16'hbd70;
mem_array[29425] = 16'h2cae;
mem_array[29424] = 16'h3e3f;
mem_array[29427] = 16'hf064;
mem_array[29426] = 16'h3ec8;
mem_array[29429] = 16'hdbdc;
mem_array[29428] = 16'hbe80;
mem_array[29431] = 16'h7a73;
mem_array[29430] = 16'h3ed1;
mem_array[29433] = 16'hff46;
mem_array[29432] = 16'hbd51;
mem_array[29435] = 16'hd48e;
mem_array[29434] = 16'h3daa;
mem_array[29437] = 16'h7390;
mem_array[29436] = 16'h3e03;
mem_array[29439] = 16'h5ab7;
mem_array[29438] = 16'h3e35;
mem_array[29441] = 16'h0cbd;
mem_array[29440] = 16'h3d03;
mem_array[29443] = 16'hec43;
mem_array[29442] = 16'h3dd2;
mem_array[29445] = 16'h9f4b;
mem_array[29444] = 16'hbcfe;
mem_array[29447] = 16'h5536;
mem_array[29446] = 16'hbd83;
mem_array[29449] = 16'h78ac;
mem_array[29448] = 16'h3e5c;
mem_array[29451] = 16'hd7e0;
mem_array[29450] = 16'h3d84;
mem_array[29453] = 16'h3d81;
mem_array[29452] = 16'hbe11;
mem_array[29455] = 16'h4734;
mem_array[29454] = 16'hbecd;
mem_array[29457] = 16'h461c;
mem_array[29456] = 16'h3e1f;
mem_array[29459] = 16'h3703;
mem_array[29458] = 16'h3e89;
mem_array[29461] = 16'hca76;
mem_array[29460] = 16'h3d9d;
mem_array[29463] = 16'hab33;
mem_array[29462] = 16'hbe71;
mem_array[29465] = 16'h1a94;
mem_array[29464] = 16'h3dc0;
mem_array[29467] = 16'h3283;
mem_array[29466] = 16'hbee6;
mem_array[29469] = 16'haa50;
mem_array[29468] = 16'h3da6;
mem_array[29471] = 16'h3478;
mem_array[29470] = 16'hbe4d;
mem_array[29473] = 16'hec50;
mem_array[29472] = 16'hbead;
mem_array[29475] = 16'hd750;
mem_array[29474] = 16'hbe41;
mem_array[29477] = 16'hab94;
mem_array[29476] = 16'h3da6;
mem_array[29479] = 16'h7373;
mem_array[29478] = 16'h3e27;
mem_array[29481] = 16'hf308;
mem_array[29480] = 16'h3d21;
mem_array[29483] = 16'h660d;
mem_array[29482] = 16'h3d08;
mem_array[29485] = 16'h31f8;
mem_array[29484] = 16'hbd83;
mem_array[29487] = 16'h14d9;
mem_array[29486] = 16'h3d68;
mem_array[29489] = 16'hc155;
mem_array[29488] = 16'hbe3d;
mem_array[29491] = 16'h668d;
mem_array[29490] = 16'h3eca;
mem_array[29493] = 16'h188b;
mem_array[29492] = 16'hbf25;
mem_array[29495] = 16'h4941;
mem_array[29494] = 16'h3d99;
mem_array[29497] = 16'hfe3d;
mem_array[29496] = 16'h3e94;
mem_array[29499] = 16'ha3cf;
mem_array[29498] = 16'h3d9f;
mem_array[29501] = 16'h8f3b;
mem_array[29500] = 16'hbd36;
mem_array[29503] = 16'h9f55;
mem_array[29502] = 16'h3e85;
mem_array[29505] = 16'haf5b;
mem_array[29504] = 16'h3e20;
mem_array[29507] = 16'hf53f;
mem_array[29506] = 16'h3c0c;
mem_array[29509] = 16'h26c8;
mem_array[29508] = 16'h3e77;
mem_array[29511] = 16'ha72a;
mem_array[29510] = 16'hbd3d;
mem_array[29513] = 16'h3382;
mem_array[29512] = 16'hbe92;
mem_array[29515] = 16'h4ab9;
mem_array[29514] = 16'h3cf0;
mem_array[29517] = 16'hc89e;
mem_array[29516] = 16'h3dda;
mem_array[29519] = 16'ha177;
mem_array[29518] = 16'h3ed8;
mem_array[29521] = 16'h862a;
mem_array[29520] = 16'hbf09;
mem_array[29523] = 16'h617d;
mem_array[29522] = 16'hbd61;
mem_array[29525] = 16'h0aa8;
mem_array[29524] = 16'h3bfe;
mem_array[29527] = 16'hfebf;
mem_array[29526] = 16'hbd37;
mem_array[29529] = 16'hff01;
mem_array[29528] = 16'hbc7c;
mem_array[29531] = 16'h42ea;
mem_array[29530] = 16'hbe23;
mem_array[29533] = 16'h3a80;
mem_array[29532] = 16'hbd07;
mem_array[29535] = 16'h2ec3;
mem_array[29534] = 16'h3d38;
mem_array[29537] = 16'h73ac;
mem_array[29536] = 16'hbddd;
mem_array[29539] = 16'hc6d4;
mem_array[29538] = 16'hbd90;
mem_array[29541] = 16'h3540;
mem_array[29540] = 16'h3cb9;
mem_array[29543] = 16'h35bb;
mem_array[29542] = 16'hbd2c;
mem_array[29545] = 16'ha126;
mem_array[29544] = 16'h3e0a;
mem_array[29547] = 16'h4e3c;
mem_array[29546] = 16'h3dd6;
mem_array[29549] = 16'h8dda;
mem_array[29548] = 16'h3e0c;
mem_array[29551] = 16'he2af;
mem_array[29550] = 16'h3e4c;
mem_array[29553] = 16'h90ec;
mem_array[29552] = 16'hbf86;
mem_array[29555] = 16'he4dc;
mem_array[29554] = 16'h3e9d;
mem_array[29557] = 16'h9cbe;
mem_array[29556] = 16'h3e20;
mem_array[29559] = 16'h22f0;
mem_array[29558] = 16'h3e12;
mem_array[29561] = 16'hee2c;
mem_array[29560] = 16'h3e86;
mem_array[29563] = 16'h06c0;
mem_array[29562] = 16'h3e21;
mem_array[29565] = 16'hc40b;
mem_array[29564] = 16'h3e98;
mem_array[29567] = 16'h3dd4;
mem_array[29566] = 16'h3dab;
mem_array[29569] = 16'hfda4;
mem_array[29568] = 16'hbb89;
mem_array[29571] = 16'hd3bf;
mem_array[29570] = 16'h3e4a;
mem_array[29573] = 16'h74f6;
mem_array[29572] = 16'hbe9b;
mem_array[29575] = 16'hbd31;
mem_array[29574] = 16'h3be2;
mem_array[29577] = 16'hd007;
mem_array[29576] = 16'h3da0;
mem_array[29579] = 16'he495;
mem_array[29578] = 16'h3e7b;
mem_array[29581] = 16'ha24e;
mem_array[29580] = 16'hbed7;
mem_array[29583] = 16'h9020;
mem_array[29582] = 16'h3caf;
mem_array[29585] = 16'hdb79;
mem_array[29584] = 16'hbe0b;
mem_array[29587] = 16'h8b71;
mem_array[29586] = 16'hbd9b;
mem_array[29589] = 16'hee4d;
mem_array[29588] = 16'h3dbb;
mem_array[29591] = 16'h1310;
mem_array[29590] = 16'h3d5f;
mem_array[29593] = 16'ha55e;
mem_array[29592] = 16'h3da3;
mem_array[29595] = 16'h2b43;
mem_array[29594] = 16'h3dad;
mem_array[29597] = 16'h37b9;
mem_array[29596] = 16'hbcd6;
mem_array[29599] = 16'hd6c5;
mem_array[29598] = 16'hbf46;
mem_array[29601] = 16'h9e82;
mem_array[29600] = 16'hbdd5;
mem_array[29603] = 16'h6e17;
mem_array[29602] = 16'hbd7f;
mem_array[29605] = 16'hc436;
mem_array[29604] = 16'h3ecb;
mem_array[29607] = 16'h255e;
mem_array[29606] = 16'hbd4b;
mem_array[29609] = 16'hbdf1;
mem_array[29608] = 16'h3db9;
mem_array[29611] = 16'ha612;
mem_array[29610] = 16'hbd37;
mem_array[29613] = 16'h0063;
mem_array[29612] = 16'hc005;
mem_array[29615] = 16'hf64c;
mem_array[29614] = 16'h3cdb;
mem_array[29617] = 16'h7994;
mem_array[29616] = 16'hbc47;
mem_array[29619] = 16'hb88e;
mem_array[29618] = 16'h3efa;
mem_array[29621] = 16'hba57;
mem_array[29620] = 16'h3e05;
mem_array[29623] = 16'h8306;
mem_array[29622] = 16'h3ed1;
mem_array[29625] = 16'hf31f;
mem_array[29624] = 16'hbd00;
mem_array[29627] = 16'hf447;
mem_array[29626] = 16'h3d62;
mem_array[29629] = 16'h0557;
mem_array[29628] = 16'hbd09;
mem_array[29631] = 16'h20dd;
mem_array[29630] = 16'hbe1e;
mem_array[29633] = 16'h7bbe;
mem_array[29632] = 16'hbe7d;
mem_array[29635] = 16'h75f3;
mem_array[29634] = 16'hbe19;
mem_array[29637] = 16'h8091;
mem_array[29636] = 16'h3d9f;
mem_array[29639] = 16'hb813;
mem_array[29638] = 16'h3e20;
mem_array[29641] = 16'h99bf;
mem_array[29640] = 16'h3eea;
mem_array[29643] = 16'hfa90;
mem_array[29642] = 16'h3d3d;
mem_array[29645] = 16'hcb3d;
mem_array[29644] = 16'h3b16;
mem_array[29647] = 16'hde87;
mem_array[29646] = 16'h3da2;
mem_array[29649] = 16'h57de;
mem_array[29648] = 16'h3d4b;
mem_array[29651] = 16'h79f9;
mem_array[29650] = 16'h3e98;
mem_array[29653] = 16'haae7;
mem_array[29652] = 16'h3e59;
mem_array[29655] = 16'h203f;
mem_array[29654] = 16'hbe2e;
mem_array[29657] = 16'hb6d1;
mem_array[29656] = 16'h3de3;
mem_array[29659] = 16'h66c9;
mem_array[29658] = 16'hbed0;
mem_array[29661] = 16'h19fe;
mem_array[29660] = 16'h3ca2;
mem_array[29663] = 16'he77d;
mem_array[29662] = 16'hbd58;
mem_array[29665] = 16'hd610;
mem_array[29664] = 16'h3ea9;
mem_array[29667] = 16'h5dd6;
mem_array[29666] = 16'h3d22;
mem_array[29669] = 16'hb0f7;
mem_array[29668] = 16'h3d31;
mem_array[29671] = 16'hbfd6;
mem_array[29670] = 16'hbdab;
mem_array[29673] = 16'hbbd7;
mem_array[29672] = 16'hbfb3;
mem_array[29675] = 16'h398e;
mem_array[29674] = 16'hbd15;
mem_array[29677] = 16'hb277;
mem_array[29676] = 16'h3e3f;
mem_array[29679] = 16'h425f;
mem_array[29678] = 16'h3e6a;
mem_array[29681] = 16'h3ff4;
mem_array[29680] = 16'hbdd4;
mem_array[29683] = 16'h4453;
mem_array[29682] = 16'h3e90;
mem_array[29685] = 16'h6289;
mem_array[29684] = 16'h3d9f;
mem_array[29687] = 16'h4498;
mem_array[29686] = 16'h3bfb;
mem_array[29689] = 16'ha401;
mem_array[29688] = 16'h3e01;
mem_array[29691] = 16'h07fd;
mem_array[29690] = 16'h3ec6;
mem_array[29693] = 16'heee3;
mem_array[29692] = 16'hbe06;
mem_array[29695] = 16'hd283;
mem_array[29694] = 16'h3e39;
mem_array[29697] = 16'he662;
mem_array[29696] = 16'h3e5b;
mem_array[29699] = 16'hf3a7;
mem_array[29698] = 16'h3e12;
mem_array[29701] = 16'haaeb;
mem_array[29700] = 16'h3e62;
mem_array[29703] = 16'h1752;
mem_array[29702] = 16'h3d96;
mem_array[29705] = 16'h8a70;
mem_array[29704] = 16'hbdac;
mem_array[29707] = 16'h2fe5;
mem_array[29706] = 16'h3dbf;
mem_array[29709] = 16'hcff1;
mem_array[29708] = 16'hbe1f;
mem_array[29711] = 16'h1d65;
mem_array[29710] = 16'h3df6;
mem_array[29713] = 16'h3b0c;
mem_array[29712] = 16'h3ecc;
mem_array[29715] = 16'h9b54;
mem_array[29714] = 16'h3db3;
mem_array[29717] = 16'ha213;
mem_array[29716] = 16'h3e91;
mem_array[29719] = 16'h591d;
mem_array[29718] = 16'h3eb7;
mem_array[29721] = 16'h23bf;
mem_array[29720] = 16'h3c9b;
mem_array[29723] = 16'hdd3f;
mem_array[29722] = 16'hbdc0;
mem_array[29725] = 16'hd64f;
mem_array[29724] = 16'h3db1;
mem_array[29727] = 16'h8ee6;
mem_array[29726] = 16'hbd57;
mem_array[29729] = 16'hd6de;
mem_array[29728] = 16'hbe49;
mem_array[29731] = 16'hed01;
mem_array[29730] = 16'hbd48;
mem_array[29733] = 16'h4da5;
mem_array[29732] = 16'hbd27;
mem_array[29735] = 16'h3546;
mem_array[29734] = 16'h3e54;
mem_array[29737] = 16'h5d96;
mem_array[29736] = 16'hbde6;
mem_array[29739] = 16'hac65;
mem_array[29738] = 16'h3ee0;
mem_array[29741] = 16'h0a70;
mem_array[29740] = 16'h3d42;
mem_array[29743] = 16'hb111;
mem_array[29742] = 16'h3f00;
mem_array[29745] = 16'h78ab;
mem_array[29744] = 16'h3ea8;
mem_array[29747] = 16'h53e7;
mem_array[29746] = 16'h3b44;
mem_array[29749] = 16'hbb9d;
mem_array[29748] = 16'hbdd8;
mem_array[29751] = 16'h7a13;
mem_array[29750] = 16'hbd04;
mem_array[29753] = 16'h1c60;
mem_array[29752] = 16'h3c05;
mem_array[29755] = 16'hbd11;
mem_array[29754] = 16'hbdb6;
mem_array[29757] = 16'hbe14;
mem_array[29756] = 16'h3e72;
mem_array[29759] = 16'hb25c;
mem_array[29758] = 16'h3eff;
mem_array[29761] = 16'h647c;
mem_array[29760] = 16'hbd95;
mem_array[29763] = 16'h050f;
mem_array[29762] = 16'h3e22;
mem_array[29765] = 16'h9246;
mem_array[29764] = 16'hbe6c;
mem_array[29767] = 16'h7ad6;
mem_array[29766] = 16'h3ea1;
mem_array[29769] = 16'he52d;
mem_array[29768] = 16'h3c9c;
mem_array[29771] = 16'h1810;
mem_array[29770] = 16'h3e89;
mem_array[29773] = 16'h82c8;
mem_array[29772] = 16'h3e28;
mem_array[29775] = 16'h7299;
mem_array[29774] = 16'hbe31;
mem_array[29777] = 16'h3055;
mem_array[29776] = 16'h3e9d;
mem_array[29779] = 16'h9603;
mem_array[29778] = 16'h3eb1;
mem_array[29781] = 16'hc6a8;
mem_array[29780] = 16'h3cd5;
mem_array[29783] = 16'h890e;
mem_array[29782] = 16'h3c56;
mem_array[29785] = 16'h3bed;
mem_array[29784] = 16'h3e8d;
mem_array[29787] = 16'h75cd;
mem_array[29786] = 16'h3e03;
mem_array[29789] = 16'hbdb4;
mem_array[29788] = 16'hbda6;
mem_array[29791] = 16'h103c;
mem_array[29790] = 16'hbd59;
mem_array[29793] = 16'h128a;
mem_array[29792] = 16'h3f09;
mem_array[29795] = 16'hd041;
mem_array[29794] = 16'hbef2;
mem_array[29797] = 16'hfe79;
mem_array[29796] = 16'hbcab;
mem_array[29799] = 16'hde30;
mem_array[29798] = 16'h3f02;
mem_array[29801] = 16'he56d;
mem_array[29800] = 16'h3f06;
mem_array[29803] = 16'h56cf;
mem_array[29802] = 16'h3f14;
mem_array[29805] = 16'h0fc2;
mem_array[29804] = 16'h3e27;
mem_array[29807] = 16'h494b;
mem_array[29806] = 16'h3e3c;
mem_array[29809] = 16'h1d28;
mem_array[29808] = 16'h3d23;
mem_array[29811] = 16'hbf2d;
mem_array[29810] = 16'hbe8c;
mem_array[29813] = 16'h2ce7;
mem_array[29812] = 16'h3d2e;
mem_array[29815] = 16'he9d7;
mem_array[29814] = 16'h3ccf;
mem_array[29817] = 16'h4c7a;
mem_array[29816] = 16'hbd2d;
mem_array[29819] = 16'h6530;
mem_array[29818] = 16'h3f06;
mem_array[29821] = 16'h66b3;
mem_array[29820] = 16'hbdeb;
mem_array[29823] = 16'h2dc6;
mem_array[29822] = 16'h3eac;
mem_array[29825] = 16'h6b29;
mem_array[29824] = 16'hbe87;
mem_array[29827] = 16'hf0de;
mem_array[29826] = 16'hbd43;
mem_array[29829] = 16'h9b04;
mem_array[29828] = 16'h3e9a;
mem_array[29831] = 16'h9283;
mem_array[29830] = 16'h3d36;
mem_array[29833] = 16'hebf4;
mem_array[29832] = 16'h3eb3;
mem_array[29835] = 16'h912c;
mem_array[29834] = 16'h3eeb;
mem_array[29837] = 16'h501d;
mem_array[29836] = 16'hbd6f;
mem_array[29839] = 16'ha585;
mem_array[29838] = 16'h3aff;
mem_array[29841] = 16'h11e0;
mem_array[29840] = 16'h3d43;
mem_array[29843] = 16'hed37;
mem_array[29842] = 16'h3d1f;
mem_array[29845] = 16'hee00;
mem_array[29844] = 16'h3e0f;
mem_array[29847] = 16'hd054;
mem_array[29846] = 16'hbe9d;
mem_array[29849] = 16'h8707;
mem_array[29848] = 16'h3ea3;
mem_array[29851] = 16'hd997;
mem_array[29850] = 16'hbe13;
mem_array[29853] = 16'had57;
mem_array[29852] = 16'h3eed;
mem_array[29855] = 16'h86a1;
mem_array[29854] = 16'h3e42;
mem_array[29857] = 16'hea55;
mem_array[29856] = 16'hbe5c;
mem_array[29859] = 16'hd06d;
mem_array[29858] = 16'h3e64;
mem_array[29861] = 16'h143a;
mem_array[29860] = 16'h3ef1;
mem_array[29863] = 16'h7b67;
mem_array[29862] = 16'h3ea3;
mem_array[29865] = 16'haa82;
mem_array[29864] = 16'h3e47;
mem_array[29867] = 16'hc57a;
mem_array[29866] = 16'h3d89;
mem_array[29869] = 16'hf5ea;
mem_array[29868] = 16'hbd99;
mem_array[29871] = 16'h3b57;
mem_array[29870] = 16'h3de5;
mem_array[29873] = 16'h2919;
mem_array[29872] = 16'hba8e;
mem_array[29875] = 16'hc3c2;
mem_array[29874] = 16'hbeea;
mem_array[29877] = 16'h0067;
mem_array[29876] = 16'h3ca2;
mem_array[29879] = 16'h8db9;
mem_array[29878] = 16'h3f12;
mem_array[29881] = 16'heb8f;
mem_array[29880] = 16'h3df3;
mem_array[29883] = 16'h9a1c;
mem_array[29882] = 16'h3e7d;
mem_array[29885] = 16'h0889;
mem_array[29884] = 16'hbea3;
mem_array[29887] = 16'h4a89;
mem_array[29886] = 16'h3d70;
mem_array[29889] = 16'h4081;
mem_array[29888] = 16'h3e2c;
mem_array[29891] = 16'h4f2b;
mem_array[29890] = 16'hbbd2;
mem_array[29893] = 16'h274e;
mem_array[29892] = 16'h3e8c;
mem_array[29895] = 16'hc757;
mem_array[29894] = 16'h3e0d;
mem_array[29897] = 16'h88fe;
mem_array[29896] = 16'hbedb;
mem_array[29899] = 16'h9dba;
mem_array[29898] = 16'hbe7b;
mem_array[29901] = 16'h8608;
mem_array[29900] = 16'h3d1d;
mem_array[29903] = 16'h5a67;
mem_array[29902] = 16'hbc3f;
mem_array[29905] = 16'h2f1a;
mem_array[29904] = 16'h3eec;
mem_array[29907] = 16'h11d8;
mem_array[29906] = 16'h3b29;
mem_array[29909] = 16'h7691;
mem_array[29908] = 16'h3e15;
mem_array[29911] = 16'hbf3c;
mem_array[29910] = 16'hbd80;
mem_array[29913] = 16'h9b75;
mem_array[29912] = 16'h3e51;
mem_array[29915] = 16'h670d;
mem_array[29914] = 16'hbe84;
mem_array[29917] = 16'h840b;
mem_array[29916] = 16'hbe10;
mem_array[29919] = 16'h4c93;
mem_array[29918] = 16'hbdc4;
mem_array[29921] = 16'hbc0f;
mem_array[29920] = 16'h3f18;
mem_array[29923] = 16'ha788;
mem_array[29922] = 16'h3e07;
mem_array[29925] = 16'h8075;
mem_array[29924] = 16'h3daf;
mem_array[29927] = 16'h7c54;
mem_array[29926] = 16'hbe25;
mem_array[29929] = 16'h1566;
mem_array[29928] = 16'hbec3;
mem_array[29931] = 16'h0eea;
mem_array[29930] = 16'hbe95;
mem_array[29933] = 16'h6f7d;
mem_array[29932] = 16'h3dcb;
mem_array[29935] = 16'he34d;
mem_array[29934] = 16'hbf90;
mem_array[29937] = 16'he08b;
mem_array[29936] = 16'h3df5;
mem_array[29939] = 16'hb30c;
mem_array[29938] = 16'h3eb8;
mem_array[29941] = 16'hcf89;
mem_array[29940] = 16'hbd3e;
mem_array[29943] = 16'hc6a3;
mem_array[29942] = 16'h3c08;
mem_array[29945] = 16'hdda1;
mem_array[29944] = 16'hbe5c;
mem_array[29947] = 16'h7072;
mem_array[29946] = 16'h3d59;
mem_array[29949] = 16'hf9cb;
mem_array[29948] = 16'h3dbd;
mem_array[29951] = 16'hc2bc;
mem_array[29950] = 16'hbdd6;
mem_array[29953] = 16'h0d08;
mem_array[29952] = 16'h3ea4;
mem_array[29955] = 16'h3420;
mem_array[29954] = 16'hbe4f;
mem_array[29957] = 16'h9b20;
mem_array[29956] = 16'h3d21;
mem_array[29959] = 16'h6904;
mem_array[29958] = 16'hbe3f;
mem_array[29961] = 16'h84db;
mem_array[29960] = 16'hbcfa;
mem_array[29963] = 16'hca89;
mem_array[29962] = 16'hbdeb;
mem_array[29965] = 16'h4111;
mem_array[29964] = 16'h3e68;
mem_array[29967] = 16'h9e5d;
mem_array[29966] = 16'h3e5b;
mem_array[29969] = 16'h33db;
mem_array[29968] = 16'h3d07;
mem_array[29971] = 16'h99d2;
mem_array[29970] = 16'h3d9c;
mem_array[29973] = 16'h0135;
mem_array[29972] = 16'h3eae;
mem_array[29975] = 16'h79ec;
mem_array[29974] = 16'hbef8;
mem_array[29977] = 16'ha7a6;
mem_array[29976] = 16'hbe88;
mem_array[29979] = 16'h1a05;
mem_array[29978] = 16'h3edc;
mem_array[29981] = 16'hff68;
mem_array[29980] = 16'h3f14;
mem_array[29983] = 16'haf73;
mem_array[29982] = 16'h3dc7;
mem_array[29985] = 16'h3a93;
mem_array[29984] = 16'hbf26;
mem_array[29987] = 16'he131;
mem_array[29986] = 16'hbe59;
mem_array[29989] = 16'hbece;
mem_array[29988] = 16'hbee8;
mem_array[29991] = 16'h818d;
mem_array[29990] = 16'hbec5;
mem_array[29993] = 16'h3df5;
mem_array[29992] = 16'hbe70;
mem_array[29995] = 16'hd4d5;
mem_array[29994] = 16'hbf8d;
mem_array[29997] = 16'h2a95;
mem_array[29996] = 16'h3edf;
mem_array[29999] = 16'h5ded;
mem_array[29998] = 16'h3eca;
mem_array[30001] = 16'h4fe9;
mem_array[30000] = 16'h3f28;
mem_array[30003] = 16'hf89a;
mem_array[30002] = 16'hbea2;
mem_array[30005] = 16'h6d5b;
mem_array[30004] = 16'h3ebb;
mem_array[30007] = 16'hedc9;
mem_array[30006] = 16'hbe11;
mem_array[30009] = 16'h2aa7;
mem_array[30008] = 16'h3e0b;
mem_array[30011] = 16'h3131;
mem_array[30010] = 16'h3f15;
mem_array[30013] = 16'hefe0;
mem_array[30012] = 16'h3e12;
mem_array[30015] = 16'h1fcb;
mem_array[30014] = 16'hbe5d;
mem_array[30017] = 16'h230f;
mem_array[30016] = 16'h3da5;
mem_array[30019] = 16'h6220;
mem_array[30018] = 16'hbf00;
mem_array[30021] = 16'h7c79;
mem_array[30020] = 16'h3c75;
mem_array[30023] = 16'hf81c;
mem_array[30022] = 16'h3cd9;
mem_array[30025] = 16'hbb78;
mem_array[30024] = 16'h3dc7;
mem_array[30027] = 16'h21a8;
mem_array[30026] = 16'h3de3;
mem_array[30029] = 16'hde1c;
mem_array[30028] = 16'hbeb3;
mem_array[30031] = 16'h3533;
mem_array[30030] = 16'h3dc6;
mem_array[30033] = 16'h53da;
mem_array[30032] = 16'hbeec;
mem_array[30035] = 16'h50a8;
mem_array[30034] = 16'hbe8f;
mem_array[30037] = 16'h34d0;
mem_array[30036] = 16'hbeed;
mem_array[30039] = 16'h1aa5;
mem_array[30038] = 16'h3e6d;
mem_array[30041] = 16'h475d;
mem_array[30040] = 16'h3ee5;
mem_array[30043] = 16'h0899;
mem_array[30042] = 16'h3e5b;
mem_array[30045] = 16'h01e0;
mem_array[30044] = 16'h3e4b;
mem_array[30047] = 16'h7fa5;
mem_array[30046] = 16'h3bb7;
mem_array[30049] = 16'h1fcf;
mem_array[30048] = 16'h3e40;
mem_array[30051] = 16'h9695;
mem_array[30050] = 16'h3d89;
mem_array[30053] = 16'h5ac2;
mem_array[30052] = 16'h3efe;
mem_array[30055] = 16'h2b4b;
mem_array[30054] = 16'hbefa;
mem_array[30057] = 16'hd32f;
mem_array[30056] = 16'h3e76;
mem_array[30059] = 16'h7875;
mem_array[30058] = 16'h3f30;
mem_array[30061] = 16'ha219;
mem_array[30060] = 16'h3f31;
mem_array[30063] = 16'h9f28;
mem_array[30062] = 16'hbf0a;
mem_array[30065] = 16'h6f62;
mem_array[30064] = 16'h3f5d;
mem_array[30067] = 16'hbe88;
mem_array[30066] = 16'hbf14;
mem_array[30069] = 16'h4971;
mem_array[30068] = 16'h3f5a;
mem_array[30071] = 16'hc079;
mem_array[30070] = 16'hbfa7;
mem_array[30073] = 16'hd376;
mem_array[30072] = 16'h3ece;
mem_array[30075] = 16'hee23;
mem_array[30074] = 16'h3f01;
mem_array[30077] = 16'h5bfa;
mem_array[30076] = 16'h3f29;
mem_array[30079] = 16'h8cd6;
mem_array[30078] = 16'hbc9e;
mem_array[30081] = 16'h9344;
mem_array[30080] = 16'hbdbb;
mem_array[30083] = 16'h2e8f;
mem_array[30082] = 16'h3c17;
mem_array[30085] = 16'h8a0d;
mem_array[30084] = 16'h3f3d;
mem_array[30087] = 16'h0f57;
mem_array[30086] = 16'h3f1e;
mem_array[30089] = 16'h0b58;
mem_array[30088] = 16'h3fab;
mem_array[30091] = 16'hc10e;
mem_array[30090] = 16'hbdd9;
mem_array[30093] = 16'h9dce;
mem_array[30092] = 16'h3ec0;
mem_array[30095] = 16'h5a64;
mem_array[30094] = 16'h3f01;
mem_array[30097] = 16'h5395;
mem_array[30096] = 16'hbf8d;
mem_array[30099] = 16'h3b59;
mem_array[30098] = 16'h3f42;
mem_array[30101] = 16'h1e1b;
mem_array[30100] = 16'h3f67;
mem_array[30103] = 16'hfa61;
mem_array[30102] = 16'hbed2;
mem_array[30105] = 16'h331f;
mem_array[30104] = 16'hbf18;
mem_array[30107] = 16'h666b;
mem_array[30106] = 16'h3dcc;
mem_array[30109] = 16'hd1eb;
mem_array[30108] = 16'h3f6a;
mem_array[30111] = 16'ha927;
mem_array[30110] = 16'h3ea3;
mem_array[30113] = 16'h61f5;
mem_array[30112] = 16'h3d86;
mem_array[30115] = 16'hc532;
mem_array[30114] = 16'hbf28;
mem_array[30117] = 16'he226;
mem_array[30116] = 16'h3f38;
mem_array[30119] = 16'h616f;
mem_array[30118] = 16'hbe43;
mem_array[30121] = 16'h739a;
mem_array[30120] = 16'h3e9e;
mem_array[30123] = 16'he9f9;
mem_array[30122] = 16'hbe1e;
mem_array[30125] = 16'h4723;
mem_array[30124] = 16'h3f59;
mem_array[30127] = 16'h2cfd;
mem_array[30126] = 16'hbfbd;
mem_array[30129] = 16'haf05;
mem_array[30128] = 16'h3f0c;
mem_array[30131] = 16'h6c88;
mem_array[30130] = 16'hbf8f;
mem_array[30133] = 16'h3f84;
mem_array[30132] = 16'h3ede;
mem_array[30135] = 16'ha5fc;
mem_array[30134] = 16'h3dfc;
mem_array[30137] = 16'hbc12;
mem_array[30136] = 16'h3f3b;
mem_array[30139] = 16'hd321;
mem_array[30138] = 16'h3ea6;
mem_array[30141] = 16'h0c0a;
mem_array[30140] = 16'hbda5;
mem_array[30143] = 16'hf598;
mem_array[30142] = 16'h3ccd;
mem_array[30145] = 16'hb183;
mem_array[30144] = 16'hbea2;
mem_array[30147] = 16'he3a6;
mem_array[30146] = 16'h3f90;
mem_array[30149] = 16'hade7;
mem_array[30148] = 16'h3f76;
mem_array[30151] = 16'hda6e;
mem_array[30150] = 16'hbe92;
mem_array[30153] = 16'ha851;
mem_array[30152] = 16'h3fa5;
mem_array[30155] = 16'h219d;
mem_array[30154] = 16'h3e03;
mem_array[30157] = 16'h918c;
mem_array[30156] = 16'hbfaf;
mem_array[30159] = 16'hc28d;
mem_array[30158] = 16'h3f46;
mem_array[30161] = 16'hb903;
mem_array[30160] = 16'h3f10;
mem_array[30163] = 16'he80e;
mem_array[30162] = 16'hbf03;
mem_array[30165] = 16'haa7c;
mem_array[30164] = 16'hbf78;
mem_array[30167] = 16'h343d;
mem_array[30166] = 16'h3e0e;
mem_array[30169] = 16'h5b0b;
mem_array[30168] = 16'h3f24;
mem_array[30171] = 16'h64fe;
mem_array[30170] = 16'h3e02;
mem_array[30173] = 16'h5314;
mem_array[30172] = 16'hbe39;
mem_array[30175] = 16'h751f;
mem_array[30174] = 16'hbef2;
mem_array[30177] = 16'h2b58;
mem_array[30176] = 16'h3f01;
mem_array[30179] = 16'hc0ed;
mem_array[30178] = 16'hbf02;
mem_array[30181] = 16'hb6bf;
mem_array[30180] = 16'h3ca5;
mem_array[30183] = 16'h0451;
mem_array[30182] = 16'h3d04;
mem_array[30185] = 16'haeef;
mem_array[30184] = 16'h3f31;
mem_array[30187] = 16'h4301;
mem_array[30186] = 16'hbf5c;
mem_array[30189] = 16'h9747;
mem_array[30188] = 16'hbdf2;
mem_array[30191] = 16'h885e;
mem_array[30190] = 16'hbe32;
mem_array[30193] = 16'h1395;
mem_array[30192] = 16'h3fc8;
mem_array[30195] = 16'h0426;
mem_array[30194] = 16'h3f24;
mem_array[30197] = 16'h387e;
mem_array[30196] = 16'h3f82;
mem_array[30199] = 16'hf224;
mem_array[30198] = 16'h3f05;
mem_array[30201] = 16'h032d;
mem_array[30200] = 16'hbd8e;
mem_array[30203] = 16'hc59c;
mem_array[30202] = 16'h3b9f;
mem_array[30205] = 16'h859a;
mem_array[30204] = 16'hbda2;
mem_array[30207] = 16'hf57c;
mem_array[30206] = 16'h3f97;
mem_array[30209] = 16'h6407;
mem_array[30208] = 16'h3e1d;
mem_array[30211] = 16'h102e;
mem_array[30210] = 16'hbf45;
mem_array[30213] = 16'h1580;
mem_array[30212] = 16'h3fc4;
mem_array[30215] = 16'h659a;
mem_array[30214] = 16'h3b18;
mem_array[30217] = 16'h851d;
mem_array[30216] = 16'hbeea;
mem_array[30219] = 16'hdbdb;
mem_array[30218] = 16'hbf1b;
mem_array[30221] = 16'h0b04;
mem_array[30220] = 16'hbe49;
mem_array[30223] = 16'hd875;
mem_array[30222] = 16'hbec7;
mem_array[30225] = 16'hcb36;
mem_array[30224] = 16'h3df1;
mem_array[30227] = 16'h630e;
mem_array[30226] = 16'hbf81;
mem_array[30229] = 16'h011a;
mem_array[30228] = 16'h3f86;
mem_array[30231] = 16'h11fe;
mem_array[30230] = 16'hbcd4;
mem_array[30233] = 16'ha06d;
mem_array[30232] = 16'h3fc7;
mem_array[30235] = 16'h6c45;
mem_array[30234] = 16'hbedd;
mem_array[30237] = 16'h0225;
mem_array[30236] = 16'h3f14;
mem_array[30239] = 16'h7308;
mem_array[30238] = 16'hbf96;
mem_array[30241] = 16'h96ce;
mem_array[30240] = 16'hbd7d;
mem_array[30243] = 16'h2701;
mem_array[30242] = 16'h3f1f;
mem_array[30245] = 16'h055e;
mem_array[30244] = 16'h3d02;
mem_array[30247] = 16'h4730;
mem_array[30246] = 16'h3cfe;
mem_array[30249] = 16'h2868;
mem_array[30248] = 16'h3d99;
mem_array[30251] = 16'hf63b;
mem_array[30250] = 16'hbb89;
mem_array[30253] = 16'h36d6;
mem_array[30252] = 16'h3f56;
mem_array[30255] = 16'h8251;
mem_array[30254] = 16'h3ece;
mem_array[30257] = 16'h07cd;
mem_array[30256] = 16'hbc8f;
mem_array[30259] = 16'hceef;
mem_array[30258] = 16'h3d22;
mem_array[30261] = 16'he8ca;
mem_array[30260] = 16'hbd3b;
mem_array[30263] = 16'h50dd;
mem_array[30262] = 16'hbcdd;
mem_array[30265] = 16'h45e9;
mem_array[30264] = 16'hbd9c;
mem_array[30267] = 16'h7db9;
mem_array[30266] = 16'hbd8f;
mem_array[30269] = 16'ha5f2;
mem_array[30268] = 16'hbcdf;
mem_array[30271] = 16'h537d;
mem_array[30270] = 16'hbf0d;
mem_array[30273] = 16'h6cca;
mem_array[30272] = 16'h3dbb;
mem_array[30275] = 16'hfd6e;
mem_array[30274] = 16'hbe17;
mem_array[30277] = 16'ha09c;
mem_array[30276] = 16'h3f4d;
mem_array[30279] = 16'h2fe1;
mem_array[30278] = 16'hbc11;
mem_array[30281] = 16'h8749;
mem_array[30280] = 16'hbf9a;
mem_array[30283] = 16'h7461;
mem_array[30282] = 16'h3f18;
mem_array[30285] = 16'hee12;
mem_array[30284] = 16'hbbc2;
mem_array[30287] = 16'h23e2;
mem_array[30286] = 16'hbf81;
mem_array[30289] = 16'hc323;
mem_array[30288] = 16'hbd93;
mem_array[30291] = 16'h6f78;
mem_array[30290] = 16'h3eb4;
mem_array[30293] = 16'hee2d;
mem_array[30292] = 16'h3f4b;
mem_array[30295] = 16'hfa27;
mem_array[30294] = 16'h3ecc;
mem_array[30297] = 16'h67a1;
mem_array[30296] = 16'hbcf1;
mem_array[30299] = 16'h820f;
mem_array[30298] = 16'hbf6a;
mem_array[30301] = 16'h04d5;
mem_array[30300] = 16'h3d02;
mem_array[30303] = 16'had84;
mem_array[30302] = 16'hbc9f;
mem_array[30305] = 16'h26a0;
mem_array[30304] = 16'hbdb0;
mem_array[30307] = 16'h7c41;
mem_array[30306] = 16'h3aca;
mem_array[30309] = 16'hbf5a;
mem_array[30308] = 16'hbd90;
mem_array[30311] = 16'h162c;
mem_array[30310] = 16'hbdb8;
mem_array[30313] = 16'h15ee;
mem_array[30312] = 16'h3f0c;
mem_array[30315] = 16'h0942;
mem_array[30314] = 16'hbe5b;
mem_array[30317] = 16'h2420;
mem_array[30316] = 16'h3b8b;
mem_array[30319] = 16'h3c18;
mem_array[30318] = 16'h3d18;
mem_array[30321] = 16'h7671;
mem_array[30320] = 16'hbc9e;
mem_array[30323] = 16'hddbe;
mem_array[30322] = 16'hbd89;
mem_array[30325] = 16'he88d;
mem_array[30324] = 16'hbe6c;
mem_array[30327] = 16'h6f35;
mem_array[30326] = 16'hbd98;
mem_array[30329] = 16'h76b7;
mem_array[30328] = 16'h3c90;
mem_array[30331] = 16'hc2e4;
mem_array[30330] = 16'hbea1;
mem_array[30333] = 16'h43c8;
mem_array[30332] = 16'h3e07;
mem_array[30335] = 16'hdd1c;
mem_array[30334] = 16'hbd86;
mem_array[30337] = 16'h2bf7;
mem_array[30336] = 16'hbe73;
mem_array[30339] = 16'h84ab;
mem_array[30338] = 16'h3d7c;
mem_array[30341] = 16'h156d;
mem_array[30340] = 16'h3d9f;
mem_array[30343] = 16'h8ee8;
mem_array[30342] = 16'h3cbb;
mem_array[30345] = 16'h0e0f;
mem_array[30344] = 16'h3c32;
mem_array[30347] = 16'h2689;
mem_array[30346] = 16'hbee5;
mem_array[30349] = 16'h4671;
mem_array[30348] = 16'h3edb;
mem_array[30351] = 16'h9095;
mem_array[30350] = 16'hbd9b;
mem_array[30353] = 16'h57d5;
mem_array[30352] = 16'h3ddd;
mem_array[30355] = 16'h8f23;
mem_array[30354] = 16'hbd9d;
mem_array[30357] = 16'he860;
mem_array[30356] = 16'h3e28;
mem_array[30359] = 16'h0174;
mem_array[30358] = 16'h3d2b;
mem_array[30361] = 16'he377;
mem_array[30360] = 16'h3d36;
mem_array[30363] = 16'h91e9;
mem_array[30362] = 16'h3ec5;
mem_array[30365] = 16'hcf85;
mem_array[30364] = 16'hbcf1;
mem_array[30367] = 16'h8b1a;
mem_array[30366] = 16'hbf31;
mem_array[30369] = 16'hc89f;
mem_array[30368] = 16'hbea6;
mem_array[30371] = 16'h7350;
mem_array[30370] = 16'hbed5;
mem_array[30373] = 16'hf13a;
mem_array[30372] = 16'hbd75;
mem_array[30375] = 16'h9f27;
mem_array[30374] = 16'hbec4;
mem_array[30377] = 16'h9f32;
mem_array[30376] = 16'hbeed;
mem_array[30379] = 16'h413b;
mem_array[30378] = 16'hbdb8;
mem_array[30381] = 16'h7d4d;
mem_array[30380] = 16'hbdce;
mem_array[30383] = 16'h1c44;
mem_array[30382] = 16'h3d80;
mem_array[30385] = 16'h1bdc;
mem_array[30384] = 16'h3dc4;
mem_array[30387] = 16'hcc08;
mem_array[30386] = 16'hbf09;
mem_array[30389] = 16'h385b;
mem_array[30388] = 16'hbb8c;
mem_array[30391] = 16'h91e7;
mem_array[30390] = 16'hbd8c;
mem_array[30393] = 16'h2284;
mem_array[30392] = 16'hbea3;
mem_array[30395] = 16'h61ab;
mem_array[30394] = 16'h3d85;
mem_array[30397] = 16'h0f33;
mem_array[30396] = 16'hbf58;
mem_array[30399] = 16'hba8b;
mem_array[30398] = 16'h3f36;
mem_array[30401] = 16'he2b1;
mem_array[30400] = 16'hbb2c;
mem_array[30403] = 16'h2d14;
mem_array[30402] = 16'hbe10;
mem_array[30405] = 16'h617e;
mem_array[30404] = 16'hbd60;
mem_array[30407] = 16'hc763;
mem_array[30406] = 16'hbed1;
mem_array[30409] = 16'h935d;
mem_array[30408] = 16'h3e99;
mem_array[30411] = 16'h260d;
mem_array[30410] = 16'h3ed8;
mem_array[30413] = 16'h7680;
mem_array[30412] = 16'hbe79;
mem_array[30415] = 16'hd048;
mem_array[30414] = 16'h3e0c;
mem_array[30417] = 16'hcd23;
mem_array[30416] = 16'hbf3d;
mem_array[30419] = 16'hac0d;
mem_array[30418] = 16'h3fbf;
mem_array[30421] = 16'hf34e;
mem_array[30420] = 16'h3f1c;
mem_array[30423] = 16'hf00c;
mem_array[30422] = 16'hbea0;
mem_array[30425] = 16'h75d3;
mem_array[30424] = 16'hbf1e;
mem_array[30427] = 16'h41af;
mem_array[30426] = 16'hbf94;
mem_array[30429] = 16'h3b7c;
mem_array[30428] = 16'h3eab;
mem_array[30431] = 16'h3577;
mem_array[30430] = 16'hbf0c;
mem_array[30433] = 16'h7278;
mem_array[30432] = 16'h3efd;
mem_array[30435] = 16'h8efb;
mem_array[30434] = 16'h3ef8;
mem_array[30437] = 16'h3626;
mem_array[30436] = 16'h3e26;
mem_array[30439] = 16'h6f07;
mem_array[30438] = 16'hbe9f;
mem_array[30441] = 16'hedc4;
mem_array[30440] = 16'h3d16;
mem_array[30443] = 16'h8bb7;
mem_array[30442] = 16'h3d70;
mem_array[30445] = 16'he4be;
mem_array[30444] = 16'hbf13;
mem_array[30447] = 16'hcb7a;
mem_array[30446] = 16'hbe43;
mem_array[30449] = 16'hf4d3;
mem_array[30448] = 16'h3e8d;
mem_array[30451] = 16'h57fd;
mem_array[30450] = 16'h3e15;
mem_array[30453] = 16'hbdcc;
mem_array[30452] = 16'hbda4;
mem_array[30455] = 16'h79c5;
mem_array[30454] = 16'h3f1e;
mem_array[30457] = 16'hfc51;
mem_array[30456] = 16'hc011;
mem_array[30459] = 16'h5d53;
mem_array[30458] = 16'h3e90;
mem_array[30461] = 16'h7cc1;
mem_array[30460] = 16'h3f6b;
mem_array[30463] = 16'h9302;
mem_array[30462] = 16'h3de8;
mem_array[30465] = 16'h364f;
mem_array[30464] = 16'hbf04;
mem_array[30467] = 16'h5902;
mem_array[30466] = 16'hbf1c;
mem_array[30469] = 16'h766b;
mem_array[30468] = 16'h3f57;
mem_array[30471] = 16'hc09c;
mem_array[30470] = 16'hbf83;
mem_array[30473] = 16'h9fe6;
mem_array[30472] = 16'h3ed6;
mem_array[30475] = 16'h54d8;
mem_array[30474] = 16'h3ea4;
mem_array[30477] = 16'h97f8;
mem_array[30476] = 16'h3e4d;
mem_array[30479] = 16'h9d57;
mem_array[30478] = 16'h3f04;
mem_array[30481] = 16'hc996;
mem_array[30480] = 16'hbeae;
mem_array[30483] = 16'h89b0;
mem_array[30482] = 16'h3eff;
mem_array[30485] = 16'h3621;
mem_array[30484] = 16'hbf02;
mem_array[30487] = 16'h44c3;
mem_array[30486] = 16'h3c94;
mem_array[30489] = 16'h4296;
mem_array[30488] = 16'h3e95;
mem_array[30491] = 16'h7619;
mem_array[30490] = 16'h3f05;
mem_array[30493] = 16'h5e3f;
mem_array[30492] = 16'hbf45;
mem_array[30495] = 16'he5c3;
mem_array[30494] = 16'hbdf7;
mem_array[30497] = 16'h0efd;
mem_array[30496] = 16'h3e8a;
mem_array[30499] = 16'hba75;
mem_array[30498] = 16'hbdeb;
mem_array[30501] = 16'h158e;
mem_array[30500] = 16'hbd0d;
mem_array[30503] = 16'hf9ec;
mem_array[30502] = 16'h3d46;
mem_array[30505] = 16'h231c;
mem_array[30504] = 16'h3ecd;
mem_array[30507] = 16'ha15c;
mem_array[30506] = 16'hbe06;
mem_array[30509] = 16'hfe55;
mem_array[30508] = 16'hbcfe;
mem_array[30511] = 16'h3b21;
mem_array[30510] = 16'hbc9d;
mem_array[30513] = 16'h896c;
mem_array[30512] = 16'h3eeb;
mem_array[30515] = 16'hf2fe;
mem_array[30514] = 16'h3e54;
mem_array[30517] = 16'h672e;
mem_array[30516] = 16'hbf21;
mem_array[30519] = 16'h4ea1;
mem_array[30518] = 16'hbd50;
mem_array[30521] = 16'h9397;
mem_array[30520] = 16'h3f0c;
mem_array[30523] = 16'h40b7;
mem_array[30522] = 16'h3d9f;
mem_array[30525] = 16'h5c7a;
mem_array[30524] = 16'hbf24;
mem_array[30527] = 16'h9e60;
mem_array[30526] = 16'h3ebb;
mem_array[30529] = 16'h95df;
mem_array[30528] = 16'h3eab;
mem_array[30531] = 16'h1616;
mem_array[30530] = 16'hbe43;
mem_array[30533] = 16'ha900;
mem_array[30532] = 16'h3edc;
mem_array[30535] = 16'h6f5b;
mem_array[30534] = 16'h3e52;
mem_array[30537] = 16'h36d2;
mem_array[30536] = 16'h3ec8;
mem_array[30539] = 16'hb3ea;
mem_array[30538] = 16'h3e82;
mem_array[30541] = 16'ha2d4;
mem_array[30540] = 16'hbf93;
mem_array[30543] = 16'h0733;
mem_array[30542] = 16'h3ea3;
mem_array[30545] = 16'h3c1d;
mem_array[30544] = 16'hbed9;
mem_array[30547] = 16'h3439;
mem_array[30546] = 16'h3e29;
mem_array[30549] = 16'hea21;
mem_array[30548] = 16'hbcea;
mem_array[30551] = 16'hf3ee;
mem_array[30550] = 16'h3e9a;
mem_array[30553] = 16'h0b93;
mem_array[30552] = 16'h3e78;
mem_array[30555] = 16'h9c13;
mem_array[30554] = 16'h3f07;
mem_array[30557] = 16'h82d1;
mem_array[30556] = 16'h3e81;
mem_array[30559] = 16'h3b1a;
mem_array[30558] = 16'h3d98;
mem_array[30561] = 16'h4086;
mem_array[30560] = 16'hbc85;
mem_array[30563] = 16'h5a9f;
mem_array[30562] = 16'h3daa;
mem_array[30565] = 16'h9b0e;
mem_array[30564] = 16'hbe20;
mem_array[30567] = 16'h9648;
mem_array[30566] = 16'hbd80;
mem_array[30569] = 16'hb9cc;
mem_array[30568] = 16'hbc8c;
mem_array[30571] = 16'ha617;
mem_array[30570] = 16'h3dbf;
mem_array[30573] = 16'h22e6;
mem_array[30572] = 16'hbf43;
mem_array[30575] = 16'h62e3;
mem_array[30574] = 16'h3d0c;
mem_array[30577] = 16'hfd02;
mem_array[30576] = 16'h3dcf;
mem_array[30579] = 16'hdc46;
mem_array[30578] = 16'h3dc0;
mem_array[30581] = 16'hdc8f;
mem_array[30580] = 16'hbe47;
mem_array[30583] = 16'h082c;
mem_array[30582] = 16'h3e84;
mem_array[30585] = 16'h52ce;
mem_array[30584] = 16'hbefa;
mem_array[30587] = 16'ha257;
mem_array[30586] = 16'h3e9e;
mem_array[30589] = 16'h8477;
mem_array[30588] = 16'h3c77;
mem_array[30591] = 16'h07ab;
mem_array[30590] = 16'hbe0f;
mem_array[30593] = 16'hc356;
mem_array[30592] = 16'h3e80;
mem_array[30595] = 16'h0ed6;
mem_array[30594] = 16'h3e5d;
mem_array[30597] = 16'h286b;
mem_array[30596] = 16'h3ed5;
mem_array[30599] = 16'h0a9e;
mem_array[30598] = 16'hbe9f;
mem_array[30601] = 16'h3bb0;
mem_array[30600] = 16'hbf4b;
mem_array[30603] = 16'hb38f;
mem_array[30602] = 16'h3e4f;
mem_array[30605] = 16'hc9ff;
mem_array[30604] = 16'hbe25;
mem_array[30607] = 16'h5414;
mem_array[30606] = 16'h3e35;
mem_array[30609] = 16'h230c;
mem_array[30608] = 16'hbdfe;
mem_array[30611] = 16'hca76;
mem_array[30610] = 16'h3e3e;
mem_array[30613] = 16'h97fd;
mem_array[30612] = 16'h3f0f;
mem_array[30615] = 16'h57b9;
mem_array[30614] = 16'h3e9b;
mem_array[30617] = 16'hfeb7;
mem_array[30616] = 16'h3e96;
mem_array[30619] = 16'haa69;
mem_array[30618] = 16'hbfac;
mem_array[30621] = 16'h293a;
mem_array[30620] = 16'hbca4;
mem_array[30623] = 16'h51c3;
mem_array[30622] = 16'h3c93;
mem_array[30625] = 16'h4675;
mem_array[30624] = 16'hbd1a;
mem_array[30627] = 16'hea5e;
mem_array[30626] = 16'h3f05;
mem_array[30629] = 16'h2518;
mem_array[30628] = 16'h3e23;
mem_array[30631] = 16'hd7e0;
mem_array[30630] = 16'h3e0b;
mem_array[30633] = 16'h746f;
mem_array[30632] = 16'hbebd;
mem_array[30635] = 16'h1419;
mem_array[30634] = 16'h3e56;
mem_array[30637] = 16'hbfc5;
mem_array[30636] = 16'h3e30;
mem_array[30639] = 16'hee32;
mem_array[30638] = 16'h3e91;
mem_array[30641] = 16'h105e;
mem_array[30640] = 16'hbccb;
mem_array[30643] = 16'hd3ee;
mem_array[30642] = 16'h3e9a;
mem_array[30645] = 16'h75ac;
mem_array[30644] = 16'hbfa1;
mem_array[30647] = 16'h6ab5;
mem_array[30646] = 16'h3e47;
mem_array[30649] = 16'h8ec2;
mem_array[30648] = 16'hbea4;
mem_array[30651] = 16'h1cd1;
mem_array[30650] = 16'hbed8;
mem_array[30653] = 16'hf73e;
mem_array[30652] = 16'h3c62;
mem_array[30655] = 16'h0b1e;
mem_array[30654] = 16'hbdab;
mem_array[30657] = 16'ha13b;
mem_array[30656] = 16'h3db9;
mem_array[30659] = 16'h7b80;
mem_array[30658] = 16'h3d9c;
mem_array[30661] = 16'hee3f;
mem_array[30660] = 16'hbeef;
mem_array[30663] = 16'h1e79;
mem_array[30662] = 16'h3e9a;
mem_array[30665] = 16'h3780;
mem_array[30664] = 16'h3f04;
mem_array[30667] = 16'h48f0;
mem_array[30666] = 16'h3e94;
mem_array[30669] = 16'h6e1c;
mem_array[30668] = 16'h3dc9;
mem_array[30671] = 16'hdd9d;
mem_array[30670] = 16'h3eed;
mem_array[30673] = 16'hbc16;
mem_array[30672] = 16'h3e83;
mem_array[30675] = 16'h78fe;
mem_array[30674] = 16'h3e90;
mem_array[30677] = 16'h0d34;
mem_array[30676] = 16'h3d74;
mem_array[30679] = 16'h9fd0;
mem_array[30678] = 16'hbea5;
mem_array[30681] = 16'h0c39;
mem_array[30680] = 16'h3cc1;
mem_array[30683] = 16'h86a4;
mem_array[30682] = 16'h3d11;
mem_array[30685] = 16'h726f;
mem_array[30684] = 16'h3eac;
mem_array[30687] = 16'h1b07;
mem_array[30686] = 16'h3ecf;
mem_array[30689] = 16'h700b;
mem_array[30688] = 16'h3e3f;
mem_array[30691] = 16'h6564;
mem_array[30690] = 16'h3e32;
mem_array[30693] = 16'h3204;
mem_array[30692] = 16'hbe95;
mem_array[30695] = 16'hef2a;
mem_array[30694] = 16'h3e51;
mem_array[30697] = 16'h95e2;
mem_array[30696] = 16'h3f0c;
mem_array[30699] = 16'h0713;
mem_array[30698] = 16'h3ed0;
mem_array[30701] = 16'h8467;
mem_array[30700] = 16'hbeae;
mem_array[30703] = 16'hfc70;
mem_array[30702] = 16'hbe14;
mem_array[30705] = 16'h5199;
mem_array[30704] = 16'hbe71;
mem_array[30707] = 16'h581a;
mem_array[30706] = 16'h3ee6;
mem_array[30709] = 16'h1065;
mem_array[30708] = 16'hbef8;
mem_array[30711] = 16'ha80a;
mem_array[30710] = 16'h3d69;
mem_array[30713] = 16'hc863;
mem_array[30712] = 16'hbeb1;
mem_array[30715] = 16'h8866;
mem_array[30714] = 16'hbee0;
mem_array[30717] = 16'ha564;
mem_array[30716] = 16'h3e1d;
mem_array[30719] = 16'h2c7b;
mem_array[30718] = 16'h3f06;
mem_array[30721] = 16'hdfe7;
mem_array[30720] = 16'hbdfa;
mem_array[30723] = 16'h9bd7;
mem_array[30722] = 16'h3ec5;
mem_array[30725] = 16'h22fb;
mem_array[30724] = 16'hbe5f;
mem_array[30727] = 16'h1893;
mem_array[30726] = 16'h3f0e;
mem_array[30729] = 16'h6468;
mem_array[30728] = 16'hbe86;
mem_array[30731] = 16'hbb12;
mem_array[30730] = 16'h3ee3;
mem_array[30733] = 16'h5d38;
mem_array[30732] = 16'h3e44;
mem_array[30735] = 16'h5b5d;
mem_array[30734] = 16'h3f02;
mem_array[30737] = 16'h4fc9;
mem_array[30736] = 16'h3d66;
mem_array[30739] = 16'h410c;
mem_array[30738] = 16'h3dde;
mem_array[30741] = 16'h5507;
mem_array[30740] = 16'hbd4e;
mem_array[30743] = 16'h8a21;
mem_array[30742] = 16'h3c51;
mem_array[30745] = 16'h782e;
mem_array[30744] = 16'h3e0b;
mem_array[30747] = 16'h0841;
mem_array[30746] = 16'h3ec6;
mem_array[30749] = 16'hacd2;
mem_array[30748] = 16'h3ebf;
mem_array[30751] = 16'hc295;
mem_array[30750] = 16'h3e82;
mem_array[30753] = 16'h910e;
mem_array[30752] = 16'h3e29;
mem_array[30755] = 16'h1c9e;
mem_array[30754] = 16'hbd60;
mem_array[30757] = 16'hca69;
mem_array[30756] = 16'h3e40;
mem_array[30759] = 16'h1588;
mem_array[30758] = 16'h3e9c;
mem_array[30761] = 16'h4970;
mem_array[30760] = 16'hbf10;
mem_array[30763] = 16'h1d32;
mem_array[30762] = 16'hbc8c;
mem_array[30765] = 16'h3f32;
mem_array[30764] = 16'hbd8a;
mem_array[30767] = 16'h812b;
mem_array[30766] = 16'h3f09;
mem_array[30769] = 16'h5a62;
mem_array[30768] = 16'hbf07;
mem_array[30771] = 16'hd9cb;
mem_array[30770] = 16'hbe4b;
mem_array[30773] = 16'hc90c;
mem_array[30772] = 16'hbe27;
mem_array[30775] = 16'h21e9;
mem_array[30774] = 16'hbf1b;
mem_array[30777] = 16'h805b;
mem_array[30776] = 16'h3e8e;
mem_array[30779] = 16'h3eb2;
mem_array[30778] = 16'h3d82;
mem_array[30781] = 16'he832;
mem_array[30780] = 16'h3d0d;
mem_array[30783] = 16'h1338;
mem_array[30782] = 16'hbe4c;
mem_array[30785] = 16'h1d76;
mem_array[30784] = 16'h3d4c;
mem_array[30787] = 16'h7eb1;
mem_array[30786] = 16'h3f2a;
mem_array[30789] = 16'h8b7a;
mem_array[30788] = 16'hbf1a;
mem_array[30791] = 16'h1465;
mem_array[30790] = 16'hbe7f;
mem_array[30793] = 16'h2a61;
mem_array[30792] = 16'h3d09;
mem_array[30795] = 16'h8bd4;
mem_array[30794] = 16'h3f12;
mem_array[30797] = 16'h4052;
mem_array[30796] = 16'hbcc6;
mem_array[30799] = 16'he9a2;
mem_array[30798] = 16'h3da6;
mem_array[30801] = 16'hf9f8;
mem_array[30800] = 16'h3c4d;
mem_array[30803] = 16'h0668;
mem_array[30802] = 16'h3d1c;
mem_array[30805] = 16'h3b24;
mem_array[30804] = 16'h3def;
mem_array[30807] = 16'h3882;
mem_array[30806] = 16'h3e51;
mem_array[30809] = 16'h2c92;
mem_array[30808] = 16'h3e97;
mem_array[30811] = 16'h0b3c;
mem_array[30810] = 16'h3f33;
mem_array[30813] = 16'hd822;
mem_array[30812] = 16'h3ea9;
mem_array[30815] = 16'h961a;
mem_array[30814] = 16'h3e45;
mem_array[30817] = 16'hcad6;
mem_array[30816] = 16'h3ea6;
mem_array[30819] = 16'hb154;
mem_array[30818] = 16'h3e9f;
mem_array[30821] = 16'h250a;
mem_array[30820] = 16'hbf08;
mem_array[30823] = 16'h6e8a;
mem_array[30822] = 16'h3e31;
mem_array[30825] = 16'ha2c9;
mem_array[30824] = 16'hbb1c;
mem_array[30827] = 16'h2917;
mem_array[30826] = 16'h3ef3;
mem_array[30829] = 16'h831c;
mem_array[30828] = 16'hbce8;
mem_array[30831] = 16'h83ac;
mem_array[30830] = 16'h3e4b;
mem_array[30833] = 16'h0ba4;
mem_array[30832] = 16'hbe24;
mem_array[30835] = 16'h151c;
mem_array[30834] = 16'hbf14;
mem_array[30837] = 16'h51cd;
mem_array[30836] = 16'h3d83;
mem_array[30839] = 16'hcb3c;
mem_array[30838] = 16'h3e96;
mem_array[30841] = 16'hdf82;
mem_array[30840] = 16'h3e21;
mem_array[30843] = 16'h8a7e;
mem_array[30842] = 16'hbf6c;
mem_array[30845] = 16'hed47;
mem_array[30844] = 16'h3e38;
mem_array[30847] = 16'h7379;
mem_array[30846] = 16'h3f13;
mem_array[30849] = 16'hc0e2;
mem_array[30848] = 16'hbe26;
mem_array[30851] = 16'h3549;
mem_array[30850] = 16'hbf1c;
mem_array[30853] = 16'h09ac;
mem_array[30852] = 16'hbe1b;
mem_array[30855] = 16'h7e64;
mem_array[30854] = 16'h3ef6;
mem_array[30857] = 16'he697;
mem_array[30856] = 16'hbe1f;
mem_array[30859] = 16'h3ec0;
mem_array[30858] = 16'hbdae;
mem_array[30861] = 16'h866a;
mem_array[30860] = 16'hbc63;
mem_array[30863] = 16'h132c;
mem_array[30862] = 16'h3cd2;
mem_array[30865] = 16'h304e;
mem_array[30864] = 16'h3ed0;
mem_array[30867] = 16'hb4bd;
mem_array[30866] = 16'h3d05;
mem_array[30869] = 16'hf965;
mem_array[30868] = 16'h3e0f;
mem_array[30871] = 16'h0e8a;
mem_array[30870] = 16'h3f5a;
mem_array[30873] = 16'h2556;
mem_array[30872] = 16'h3eb0;
mem_array[30875] = 16'hb8f3;
mem_array[30874] = 16'hbd6b;
mem_array[30877] = 16'hd735;
mem_array[30876] = 16'h3ec1;
mem_array[30879] = 16'hdf3e;
mem_array[30878] = 16'hbe3b;
mem_array[30881] = 16'h1e96;
mem_array[30880] = 16'hbe54;
mem_array[30883] = 16'he71a;
mem_array[30882] = 16'h3e9b;
mem_array[30885] = 16'ha3c1;
mem_array[30884] = 16'h3e55;
mem_array[30887] = 16'h9a2f;
mem_array[30886] = 16'h3f01;
mem_array[30889] = 16'hcb45;
mem_array[30888] = 16'hbef6;
mem_array[30891] = 16'h4739;
mem_array[30890] = 16'h3ed9;
mem_array[30893] = 16'h8756;
mem_array[30892] = 16'hbddb;
mem_array[30895] = 16'h5ad6;
mem_array[30894] = 16'hbec8;
mem_array[30897] = 16'hc4f0;
mem_array[30896] = 16'hbe20;
mem_array[30899] = 16'hfee6;
mem_array[30898] = 16'h3efd;
mem_array[30901] = 16'hb1ee;
mem_array[30900] = 16'h3ec5;
mem_array[30903] = 16'ha046;
mem_array[30902] = 16'hbfa7;
mem_array[30905] = 16'h5511;
mem_array[30904] = 16'h3ed3;
mem_array[30907] = 16'he22e;
mem_array[30906] = 16'hbd34;
mem_array[30909] = 16'h8798;
mem_array[30908] = 16'hbe89;
mem_array[30911] = 16'h9363;
mem_array[30910] = 16'hbf05;
mem_array[30913] = 16'hb75d;
mem_array[30912] = 16'h3c26;
mem_array[30915] = 16'h20f3;
mem_array[30914] = 16'h3eff;
mem_array[30917] = 16'h51d7;
mem_array[30916] = 16'hbd7c;
mem_array[30919] = 16'h4acc;
mem_array[30918] = 16'hbe4c;
mem_array[30921] = 16'hb29e;
mem_array[30920] = 16'hbd7a;
mem_array[30923] = 16'h165d;
mem_array[30922] = 16'hbdb1;
mem_array[30925] = 16'h5e4d;
mem_array[30924] = 16'h3eaf;
mem_array[30927] = 16'h6e26;
mem_array[30926] = 16'h3e82;
mem_array[30929] = 16'hf205;
mem_array[30928] = 16'h3e58;
mem_array[30931] = 16'ha35e;
mem_array[30930] = 16'h3f57;
mem_array[30933] = 16'h7af9;
mem_array[30932] = 16'h3f13;
mem_array[30935] = 16'hc4cc;
mem_array[30934] = 16'hbe1c;
mem_array[30937] = 16'hd20a;
mem_array[30936] = 16'h3dd8;
mem_array[30939] = 16'h6eed;
mem_array[30938] = 16'hbe8c;
mem_array[30941] = 16'ha5c5;
mem_array[30940] = 16'hbc2f;
mem_array[30943] = 16'h49e0;
mem_array[30942] = 16'h3e68;
mem_array[30945] = 16'hfea9;
mem_array[30944] = 16'h3ed2;
mem_array[30947] = 16'h25bd;
mem_array[30946] = 16'h3f2b;
mem_array[30949] = 16'h78c9;
mem_array[30948] = 16'hbed0;
mem_array[30951] = 16'h35f4;
mem_array[30950] = 16'hbe02;
mem_array[30953] = 16'h91e5;
mem_array[30952] = 16'h3dc1;
mem_array[30955] = 16'h36cb;
mem_array[30954] = 16'hbe6f;
mem_array[30957] = 16'h8e18;
mem_array[30956] = 16'hbe4f;
mem_array[30959] = 16'hdbbb;
mem_array[30958] = 16'h3e08;
mem_array[30961] = 16'hf044;
mem_array[30960] = 16'h3ec7;
mem_array[30963] = 16'hec54;
mem_array[30962] = 16'hbf03;
mem_array[30965] = 16'hc184;
mem_array[30964] = 16'h3ea6;
mem_array[30967] = 16'h5c3f;
mem_array[30966] = 16'hbf4f;
mem_array[30969] = 16'hbd6e;
mem_array[30968] = 16'h3e8c;
mem_array[30971] = 16'h5e61;
mem_array[30970] = 16'hbf34;
mem_array[30973] = 16'h6091;
mem_array[30972] = 16'hbe70;
mem_array[30975] = 16'h140a;
mem_array[30974] = 16'h3f34;
mem_array[30977] = 16'hb9cc;
mem_array[30976] = 16'hbc82;
mem_array[30979] = 16'h3bfd;
mem_array[30978] = 16'hbe84;
mem_array[30981] = 16'ha13d;
mem_array[30980] = 16'hbc3f;
mem_array[30983] = 16'h4b36;
mem_array[30982] = 16'hbbe1;
mem_array[30985] = 16'hc645;
mem_array[30984] = 16'hbd7f;
mem_array[30987] = 16'h990b;
mem_array[30986] = 16'h3e8b;
mem_array[30989] = 16'h4174;
mem_array[30988] = 16'h3e85;
mem_array[30991] = 16'h4fec;
mem_array[30990] = 16'h3f49;
mem_array[30993] = 16'h5a88;
mem_array[30992] = 16'h3e5d;
mem_array[30995] = 16'hfd22;
mem_array[30994] = 16'hbd8a;
mem_array[30997] = 16'h91c9;
mem_array[30996] = 16'hbe2d;
mem_array[30999] = 16'h6205;
mem_array[30998] = 16'hbe09;
mem_array[31001] = 16'h01f6;
mem_array[31000] = 16'h3db7;
mem_array[31003] = 16'h8adb;
mem_array[31002] = 16'h3ebb;
mem_array[31005] = 16'hf07e;
mem_array[31004] = 16'h3f10;
mem_array[31007] = 16'h84fd;
mem_array[31006] = 16'h3f29;
mem_array[31009] = 16'h72ba;
mem_array[31008] = 16'hbdc2;
mem_array[31011] = 16'h4105;
mem_array[31010] = 16'hbe89;
mem_array[31013] = 16'h2f50;
mem_array[31012] = 16'h3e3f;
mem_array[31015] = 16'h9867;
mem_array[31014] = 16'h3e6d;
mem_array[31017] = 16'h456a;
mem_array[31016] = 16'hbe0b;
mem_array[31019] = 16'h3dac;
mem_array[31018] = 16'h3eee;
mem_array[31021] = 16'h9856;
mem_array[31020] = 16'h3e6e;
mem_array[31023] = 16'h0175;
mem_array[31022] = 16'h3edb;
mem_array[31025] = 16'ha551;
mem_array[31024] = 16'h3ec6;
mem_array[31027] = 16'h19e0;
mem_array[31026] = 16'hbf12;
mem_array[31029] = 16'h0f92;
mem_array[31028] = 16'h3eb2;
mem_array[31031] = 16'h3dfd;
mem_array[31030] = 16'hbe25;
mem_array[31033] = 16'h7158;
mem_array[31032] = 16'hbf19;
mem_array[31035] = 16'h1913;
mem_array[31034] = 16'h3ed9;
mem_array[31037] = 16'h25f0;
mem_array[31036] = 16'hbe99;
mem_array[31039] = 16'hf0a1;
mem_array[31038] = 16'h3e92;
mem_array[31041] = 16'h0053;
mem_array[31040] = 16'hbd72;
mem_array[31043] = 16'h65eb;
mem_array[31042] = 16'hbd95;
mem_array[31045] = 16'hc8b5;
mem_array[31044] = 16'h3e7f;
mem_array[31047] = 16'h50d9;
mem_array[31046] = 16'h3e9e;
mem_array[31049] = 16'h3c5f;
mem_array[31048] = 16'hbc3a;
mem_array[31051] = 16'ha5ca;
mem_array[31050] = 16'h3f28;
mem_array[31053] = 16'h7843;
mem_array[31052] = 16'hbe57;
mem_array[31055] = 16'hd12a;
mem_array[31054] = 16'h3e82;
mem_array[31057] = 16'ha709;
mem_array[31056] = 16'h3e84;
mem_array[31059] = 16'he28b;
mem_array[31058] = 16'h3e02;
mem_array[31061] = 16'h1538;
mem_array[31060] = 16'h3d69;
mem_array[31063] = 16'hd0a6;
mem_array[31062] = 16'h3e90;
mem_array[31065] = 16'hf6a1;
mem_array[31064] = 16'hbe9b;
mem_array[31067] = 16'h0fbc;
mem_array[31066] = 16'h3e86;
mem_array[31069] = 16'h4d7a;
mem_array[31068] = 16'hbe16;
mem_array[31071] = 16'h6ef3;
mem_array[31070] = 16'h3eaf;
mem_array[31073] = 16'h7f5b;
mem_array[31072] = 16'h3d02;
mem_array[31075] = 16'ha710;
mem_array[31074] = 16'h3d63;
mem_array[31077] = 16'h66b3;
mem_array[31076] = 16'hbda6;
mem_array[31079] = 16'h5597;
mem_array[31078] = 16'h3f22;
mem_array[31081] = 16'h8658;
mem_array[31080] = 16'h3c00;
mem_array[31083] = 16'h6e97;
mem_array[31082] = 16'h3ef0;
mem_array[31085] = 16'hb76c;
mem_array[31084] = 16'h3e9d;
mem_array[31087] = 16'hd2d0;
mem_array[31086] = 16'hbec7;
mem_array[31089] = 16'hb144;
mem_array[31088] = 16'hbe16;
mem_array[31091] = 16'h4858;
mem_array[31090] = 16'hbce0;
mem_array[31093] = 16'h298e;
mem_array[31092] = 16'hbf1d;
mem_array[31095] = 16'ha3bb;
mem_array[31094] = 16'h3e2d;
mem_array[31097] = 16'hd005;
mem_array[31096] = 16'hbd96;
mem_array[31099] = 16'h6b17;
mem_array[31098] = 16'h3ee0;
mem_array[31101] = 16'hb7d1;
mem_array[31100] = 16'hbe37;
mem_array[31103] = 16'hb5f1;
mem_array[31102] = 16'h3ce5;
mem_array[31105] = 16'hd60c;
mem_array[31104] = 16'h3efa;
mem_array[31107] = 16'hcc8d;
mem_array[31106] = 16'h3e78;
mem_array[31109] = 16'h0c3a;
mem_array[31108] = 16'h3d5f;
mem_array[31111] = 16'h465f;
mem_array[31110] = 16'h3e9d;
mem_array[31113] = 16'h4b1c;
mem_array[31112] = 16'h3d15;
mem_array[31115] = 16'h343c;
mem_array[31114] = 16'h3e17;
mem_array[31117] = 16'h9105;
mem_array[31116] = 16'h3eaf;
mem_array[31119] = 16'hcdb8;
mem_array[31118] = 16'h3d83;
mem_array[31121] = 16'h9cb8;
mem_array[31120] = 16'hbe48;
mem_array[31123] = 16'he7da;
mem_array[31122] = 16'h3db2;
mem_array[31125] = 16'hd24a;
mem_array[31124] = 16'h3e9c;
mem_array[31127] = 16'hfa64;
mem_array[31126] = 16'h3ee8;
mem_array[31129] = 16'h7292;
mem_array[31128] = 16'hbdb0;
mem_array[31131] = 16'h1b14;
mem_array[31130] = 16'h3eda;
mem_array[31133] = 16'h1aaa;
mem_array[31132] = 16'hbeb4;
mem_array[31135] = 16'hb8b1;
mem_array[31134] = 16'hbdd7;
mem_array[31137] = 16'h13c4;
mem_array[31136] = 16'hbd84;
mem_array[31139] = 16'h37ee;
mem_array[31138] = 16'h3e21;
mem_array[31141] = 16'h376b;
mem_array[31140] = 16'hbee6;
mem_array[31143] = 16'hfd75;
mem_array[31142] = 16'hbe12;
mem_array[31145] = 16'hb43b;
mem_array[31144] = 16'h3e1e;
mem_array[31147] = 16'hfc17;
mem_array[31146] = 16'h3bbb;
mem_array[31149] = 16'h46af;
mem_array[31148] = 16'hbdd0;
mem_array[31151] = 16'hef24;
mem_array[31150] = 16'h3d66;
mem_array[31153] = 16'hf730;
mem_array[31152] = 16'hbe3a;
mem_array[31155] = 16'h78c6;
mem_array[31154] = 16'h3d35;
mem_array[31157] = 16'h8ea9;
mem_array[31156] = 16'h3c79;
mem_array[31159] = 16'hd2ee;
mem_array[31158] = 16'h3d62;
mem_array[31161] = 16'ha6c0;
mem_array[31160] = 16'hbdf8;
mem_array[31163] = 16'h0547;
mem_array[31162] = 16'hbd85;
mem_array[31165] = 16'hfe76;
mem_array[31164] = 16'h3e59;
mem_array[31167] = 16'h39ee;
mem_array[31166] = 16'h3dc3;
mem_array[31169] = 16'hab61;
mem_array[31168] = 16'hbc0c;
mem_array[31171] = 16'h6b80;
mem_array[31170] = 16'h3eb6;
mem_array[31173] = 16'h943f;
mem_array[31172] = 16'hbf80;
mem_array[31175] = 16'h767f;
mem_array[31174] = 16'h3c98;
mem_array[31177] = 16'he8b7;
mem_array[31176] = 16'h3e1f;
mem_array[31179] = 16'hf9c5;
mem_array[31178] = 16'hbcfe;
mem_array[31181] = 16'h215f;
mem_array[31180] = 16'hbd01;
mem_array[31183] = 16'hd224;
mem_array[31182] = 16'h3e6b;
mem_array[31185] = 16'h1a02;
mem_array[31184] = 16'h3ea8;
mem_array[31187] = 16'ha939;
mem_array[31186] = 16'h3ea9;
mem_array[31189] = 16'h3798;
mem_array[31188] = 16'h3e0d;
mem_array[31191] = 16'h1d08;
mem_array[31190] = 16'hbe67;
mem_array[31193] = 16'hcd38;
mem_array[31192] = 16'hbe72;
mem_array[31195] = 16'h1b32;
mem_array[31194] = 16'hbba7;
mem_array[31197] = 16'h224c;
mem_array[31196] = 16'hbd90;
mem_array[31199] = 16'hd619;
mem_array[31198] = 16'h3dfa;
mem_array[31201] = 16'h60ab;
mem_array[31200] = 16'hbf30;
mem_array[31203] = 16'hf14b;
mem_array[31202] = 16'h3bf2;
mem_array[31205] = 16'h88b0;
mem_array[31204] = 16'h3e04;
mem_array[31207] = 16'hd331;
mem_array[31206] = 16'hbcfb;
mem_array[31209] = 16'h78c1;
mem_array[31208] = 16'h3e73;
mem_array[31211] = 16'h80ca;
mem_array[31210] = 16'h3dc0;
mem_array[31213] = 16'h0a01;
mem_array[31212] = 16'h3e28;
mem_array[31215] = 16'h433c;
mem_array[31214] = 16'h3cc5;
mem_array[31217] = 16'h269e;
mem_array[31216] = 16'hbe62;
mem_array[31219] = 16'h61b4;
mem_array[31218] = 16'hbebb;
mem_array[31221] = 16'h9406;
mem_array[31220] = 16'hbd9f;
mem_array[31223] = 16'h1d70;
mem_array[31222] = 16'hbd87;
mem_array[31225] = 16'he0b9;
mem_array[31224] = 16'h3e1d;
mem_array[31227] = 16'hdb18;
mem_array[31226] = 16'h3e4b;
mem_array[31229] = 16'hd649;
mem_array[31228] = 16'hbd5a;
mem_array[31231] = 16'ha9ce;
mem_array[31230] = 16'h3d1c;
mem_array[31233] = 16'h7823;
mem_array[31232] = 16'hbf8f;
mem_array[31235] = 16'h750a;
mem_array[31234] = 16'hbe23;
mem_array[31237] = 16'hfe34;
mem_array[31236] = 16'h3d7d;
mem_array[31239] = 16'h512d;
mem_array[31238] = 16'h3e14;
mem_array[31241] = 16'h5a02;
mem_array[31240] = 16'hbe4c;
mem_array[31243] = 16'h8248;
mem_array[31242] = 16'h3e91;
mem_array[31245] = 16'hcb4b;
mem_array[31244] = 16'h3ec3;
mem_array[31247] = 16'h8171;
mem_array[31246] = 16'hbc35;
mem_array[31249] = 16'hfdfe;
mem_array[31248] = 16'h3e66;
mem_array[31251] = 16'h3743;
mem_array[31250] = 16'h39d1;
mem_array[31253] = 16'hc8ef;
mem_array[31252] = 16'hbdfd;
mem_array[31255] = 16'h3719;
mem_array[31254] = 16'h3e01;
mem_array[31257] = 16'hfbda;
mem_array[31256] = 16'hbd41;
mem_array[31259] = 16'h1573;
mem_array[31258] = 16'hbcb0;
mem_array[31261] = 16'h36f5;
mem_array[31260] = 16'hbf02;
mem_array[31263] = 16'h7ee4;
mem_array[31262] = 16'h3d2f;
mem_array[31265] = 16'h9644;
mem_array[31264] = 16'h3d81;
mem_array[31267] = 16'h629c;
mem_array[31266] = 16'h3e39;
mem_array[31269] = 16'hbe52;
mem_array[31268] = 16'hbe73;
mem_array[31271] = 16'h3958;
mem_array[31270] = 16'h3dde;
mem_array[31273] = 16'h7127;
mem_array[31272] = 16'h3e57;
mem_array[31275] = 16'had20;
mem_array[31274] = 16'hbe03;
mem_array[31277] = 16'hb823;
mem_array[31276] = 16'hbd16;
mem_array[31279] = 16'h5637;
mem_array[31278] = 16'hbe23;
mem_array[31281] = 16'hdca6;
mem_array[31280] = 16'hbc27;
mem_array[31283] = 16'hddcf;
mem_array[31282] = 16'hbd5d;
mem_array[31285] = 16'h6729;
mem_array[31284] = 16'h3edf;
mem_array[31287] = 16'h9e7c;
mem_array[31286] = 16'hbb6f;
mem_array[31289] = 16'h3920;
mem_array[31288] = 16'hbde8;
mem_array[31291] = 16'hb75f;
mem_array[31290] = 16'hbc70;
mem_array[31293] = 16'h31c0;
mem_array[31292] = 16'hbf57;
mem_array[31295] = 16'h64a5;
mem_array[31294] = 16'hbddc;
mem_array[31297] = 16'hc853;
mem_array[31296] = 16'h3e03;
mem_array[31299] = 16'h5ffb;
mem_array[31298] = 16'h3e0e;
mem_array[31301] = 16'h27a2;
mem_array[31300] = 16'hbf0c;
mem_array[31303] = 16'hc780;
mem_array[31302] = 16'h3de9;
mem_array[31305] = 16'hf3d3;
mem_array[31304] = 16'hbe7d;
mem_array[31307] = 16'hbe84;
mem_array[31306] = 16'h3e2c;
mem_array[31309] = 16'h5158;
mem_array[31308] = 16'h3e8d;
mem_array[31311] = 16'hc32f;
mem_array[31310] = 16'hbd99;
mem_array[31313] = 16'h756e;
mem_array[31312] = 16'hbe30;
mem_array[31315] = 16'h56ba;
mem_array[31314] = 16'h3ee3;
mem_array[31317] = 16'hadd2;
mem_array[31316] = 16'hbda8;
mem_array[31319] = 16'h300d;
mem_array[31318] = 16'h3dbc;
mem_array[31321] = 16'h75cc;
mem_array[31320] = 16'h3eab;
mem_array[31323] = 16'h9cd0;
mem_array[31322] = 16'h3e5a;
mem_array[31325] = 16'h32ee;
mem_array[31324] = 16'h3e07;
mem_array[31327] = 16'h447a;
mem_array[31326] = 16'h3e42;
mem_array[31329] = 16'hc9b5;
mem_array[31328] = 16'hbe46;
mem_array[31331] = 16'h6f53;
mem_array[31330] = 16'hbdfb;
mem_array[31333] = 16'h9471;
mem_array[31332] = 16'h3e35;
mem_array[31335] = 16'he803;
mem_array[31334] = 16'hbe8e;
mem_array[31337] = 16'hd2c3;
mem_array[31336] = 16'hbd88;
mem_array[31339] = 16'h02ea;
mem_array[31338] = 16'h3e8a;
mem_array[31341] = 16'h6309;
mem_array[31340] = 16'hbbb3;
mem_array[31343] = 16'h8a83;
mem_array[31342] = 16'hbcf6;
mem_array[31345] = 16'h8051;
mem_array[31344] = 16'h3e7f;
mem_array[31347] = 16'he866;
mem_array[31346] = 16'h3df6;
mem_array[31349] = 16'hdfd7;
mem_array[31348] = 16'h3e3d;
mem_array[31351] = 16'hb6d2;
mem_array[31350] = 16'hbc7c;
mem_array[31353] = 16'hd212;
mem_array[31352] = 16'h3da9;
mem_array[31355] = 16'he84e;
mem_array[31354] = 16'h3e01;
mem_array[31357] = 16'h3002;
mem_array[31356] = 16'h3d08;
mem_array[31359] = 16'h132b;
mem_array[31358] = 16'h3e8c;
mem_array[31361] = 16'hec38;
mem_array[31360] = 16'hbe4a;
mem_array[31363] = 16'he31b;
mem_array[31362] = 16'h3de2;
mem_array[31365] = 16'haeff;
mem_array[31364] = 16'h3cb8;
mem_array[31367] = 16'h6b43;
mem_array[31366] = 16'h3ea1;
mem_array[31369] = 16'h1edf;
mem_array[31368] = 16'h3e2a;
mem_array[31371] = 16'ha2b1;
mem_array[31370] = 16'hbd89;
mem_array[31373] = 16'h2323;
mem_array[31372] = 16'h3d74;
mem_array[31375] = 16'h4b83;
mem_array[31374] = 16'h3ea0;
mem_array[31377] = 16'h4041;
mem_array[31376] = 16'h3d79;
mem_array[31379] = 16'hd24b;
mem_array[31378] = 16'h3e43;
mem_array[31381] = 16'hdb86;
mem_array[31380] = 16'hbc38;
mem_array[31383] = 16'h02e9;
mem_array[31382] = 16'hbc69;
mem_array[31385] = 16'hede7;
mem_array[31384] = 16'h3e45;
mem_array[31387] = 16'h0502;
mem_array[31386] = 16'h3e08;
mem_array[31389] = 16'hd063;
mem_array[31388] = 16'hbebe;
mem_array[31391] = 16'h3850;
mem_array[31390] = 16'hbdf2;
mem_array[31393] = 16'h917b;
mem_array[31392] = 16'h3ebd;
mem_array[31395] = 16'h9f38;
mem_array[31394] = 16'hbe31;
mem_array[31397] = 16'hcb99;
mem_array[31396] = 16'h3db4;
mem_array[31399] = 16'h7879;
mem_array[31398] = 16'hbd8d;
mem_array[31401] = 16'h7b1f;
mem_array[31400] = 16'h3d22;
mem_array[31403] = 16'ha9f2;
mem_array[31402] = 16'hbd3e;
mem_array[31405] = 16'h1d6e;
mem_array[31404] = 16'hbde7;
mem_array[31407] = 16'hff0b;
mem_array[31406] = 16'h3df1;
mem_array[31409] = 16'h52f6;
mem_array[31408] = 16'hbe21;
mem_array[31411] = 16'h777a;
mem_array[31410] = 16'hbd8d;
mem_array[31413] = 16'he9a0;
mem_array[31412] = 16'h3f17;
mem_array[31415] = 16'heb73;
mem_array[31414] = 16'h3d12;
mem_array[31417] = 16'h169b;
mem_array[31416] = 16'hbde4;
mem_array[31419] = 16'hbef1;
mem_array[31418] = 16'h3dfe;
mem_array[31421] = 16'h82e0;
mem_array[31420] = 16'hbf08;
mem_array[31423] = 16'h081c;
mem_array[31422] = 16'h3eb7;
mem_array[31425] = 16'h6aca;
mem_array[31424] = 16'h3ee8;
mem_array[31427] = 16'h167d;
mem_array[31426] = 16'h3e9f;
mem_array[31429] = 16'hf159;
mem_array[31428] = 16'h3e7d;
mem_array[31431] = 16'h076e;
mem_array[31430] = 16'hbeca;
mem_array[31433] = 16'h7d2e;
mem_array[31432] = 16'h3e1d;
mem_array[31435] = 16'hb4d2;
mem_array[31434] = 16'hbe5e;
mem_array[31437] = 16'h4ab9;
mem_array[31436] = 16'h3e33;
mem_array[31439] = 16'hd70b;
mem_array[31438] = 16'h3e89;
mem_array[31441] = 16'h2188;
mem_array[31440] = 16'hbfca;
mem_array[31443] = 16'he770;
mem_array[31442] = 16'h3ece;
mem_array[31445] = 16'h9ad5;
mem_array[31444] = 16'h3cb0;
mem_array[31447] = 16'hc39c;
mem_array[31446] = 16'h3dba;
mem_array[31449] = 16'hed13;
mem_array[31448] = 16'hbeb8;
mem_array[31451] = 16'hec52;
mem_array[31450] = 16'h3d89;
mem_array[31453] = 16'h7fda;
mem_array[31452] = 16'h3e9d;
mem_array[31455] = 16'hd4fa;
mem_array[31454] = 16'hbe1c;
mem_array[31457] = 16'hf657;
mem_array[31456] = 16'hbe28;
mem_array[31459] = 16'h2ccb;
mem_array[31458] = 16'h3ebc;
mem_array[31461] = 16'h04f2;
mem_array[31460] = 16'hbd0d;
mem_array[31463] = 16'h6997;
mem_array[31462] = 16'h3c3f;
mem_array[31465] = 16'h43ea;
mem_array[31464] = 16'hbdb1;
mem_array[31467] = 16'h0bb0;
mem_array[31466] = 16'hbe25;
mem_array[31469] = 16'h033a;
mem_array[31468] = 16'hbe85;
mem_array[31471] = 16'h06a8;
mem_array[31470] = 16'hbd76;
mem_array[31473] = 16'h4e71;
mem_array[31472] = 16'h3ee7;
mem_array[31475] = 16'heb60;
mem_array[31474] = 16'hbd3d;
mem_array[31477] = 16'hb7b9;
mem_array[31476] = 16'h3925;
mem_array[31479] = 16'h79c3;
mem_array[31478] = 16'h3d5b;
mem_array[31481] = 16'h7a9f;
mem_array[31480] = 16'hbef2;
mem_array[31483] = 16'h9425;
mem_array[31482] = 16'h3ec8;
mem_array[31485] = 16'h1ce3;
mem_array[31484] = 16'h3e49;
mem_array[31487] = 16'h1b19;
mem_array[31486] = 16'h3d8f;
mem_array[31489] = 16'he263;
mem_array[31488] = 16'hbd92;
mem_array[31491] = 16'ha63d;
mem_array[31490] = 16'h3e7a;
mem_array[31493] = 16'h32ef;
mem_array[31492] = 16'h3e9b;
mem_array[31495] = 16'h2553;
mem_array[31494] = 16'hbcae;
mem_array[31497] = 16'hdf42;
mem_array[31496] = 16'hbe39;
mem_array[31499] = 16'h324c;
mem_array[31498] = 16'h3dae;
mem_array[31501] = 16'h6810;
mem_array[31500] = 16'hbe58;
mem_array[31503] = 16'h4852;
mem_array[31502] = 16'h3f29;
mem_array[31505] = 16'h0a7c;
mem_array[31504] = 16'h3e54;
mem_array[31507] = 16'hf6ea;
mem_array[31506] = 16'h3e37;
mem_array[31509] = 16'h751e;
mem_array[31508] = 16'h3e54;
mem_array[31511] = 16'h1da6;
mem_array[31510] = 16'h3e05;
mem_array[31513] = 16'h80f1;
mem_array[31512] = 16'h3f71;
mem_array[31515] = 16'h7949;
mem_array[31514] = 16'hbe9a;
mem_array[31517] = 16'h666a;
mem_array[31516] = 16'h3db1;
mem_array[31519] = 16'h4814;
mem_array[31518] = 16'h3e82;
mem_array[31521] = 16'h42dc;
mem_array[31520] = 16'h3c4d;
mem_array[31523] = 16'hf2b2;
mem_array[31522] = 16'h3c0f;
mem_array[31525] = 16'h3a08;
mem_array[31524] = 16'hbd2d;
mem_array[31527] = 16'h7480;
mem_array[31526] = 16'hbd8e;
mem_array[31529] = 16'h165c;
mem_array[31528] = 16'h3e4c;
mem_array[31531] = 16'ha8d7;
mem_array[31530] = 16'hbdd6;
mem_array[31533] = 16'hc633;
mem_array[31532] = 16'h3f1f;
mem_array[31535] = 16'h574d;
mem_array[31534] = 16'hbd1f;
mem_array[31537] = 16'h89b2;
mem_array[31536] = 16'h3dea;
mem_array[31539] = 16'h7141;
mem_array[31538] = 16'h3e9c;
mem_array[31541] = 16'he72c;
mem_array[31540] = 16'hbeb4;
mem_array[31543] = 16'hb38f;
mem_array[31542] = 16'h3e2e;
mem_array[31545] = 16'h338e;
mem_array[31544] = 16'h3e3e;
mem_array[31547] = 16'h4ed3;
mem_array[31546] = 16'hbdb2;
mem_array[31549] = 16'h08e2;
mem_array[31548] = 16'h3d9c;
mem_array[31551] = 16'h4919;
mem_array[31550] = 16'hbea7;
mem_array[31553] = 16'hb36d;
mem_array[31552] = 16'h3dc1;
mem_array[31555] = 16'h8675;
mem_array[31554] = 16'hbe86;
mem_array[31557] = 16'hc7f3;
mem_array[31556] = 16'hb987;
mem_array[31559] = 16'h8796;
mem_array[31558] = 16'h3e86;
mem_array[31561] = 16'hf0aa;
mem_array[31560] = 16'hbf56;
mem_array[31563] = 16'h72e6;
mem_array[31562] = 16'h3f0f;
mem_array[31565] = 16'h2443;
mem_array[31564] = 16'h3d76;
mem_array[31567] = 16'h65b7;
mem_array[31566] = 16'h3e42;
mem_array[31569] = 16'hd30c;
mem_array[31568] = 16'h3dc4;
mem_array[31571] = 16'h4054;
mem_array[31570] = 16'h3d94;
mem_array[31573] = 16'h2f7e;
mem_array[31572] = 16'h3efd;
mem_array[31575] = 16'h611e;
mem_array[31574] = 16'hbe97;
mem_array[31577] = 16'h8370;
mem_array[31576] = 16'h3e22;
mem_array[31579] = 16'h1ed3;
mem_array[31578] = 16'h3eab;
mem_array[31581] = 16'ha9a3;
mem_array[31580] = 16'hbd36;
mem_array[31583] = 16'h170b;
mem_array[31582] = 16'h3ca8;
mem_array[31585] = 16'h1c6a;
mem_array[31584] = 16'hbe30;
mem_array[31587] = 16'h1202;
mem_array[31586] = 16'hbd34;
mem_array[31589] = 16'haf74;
mem_array[31588] = 16'h3d9d;
mem_array[31591] = 16'hd783;
mem_array[31590] = 16'h3dcd;
mem_array[31593] = 16'hbecb;
mem_array[31592] = 16'h3f35;
mem_array[31595] = 16'h692b;
mem_array[31594] = 16'hbf09;
mem_array[31597] = 16'he3ba;
mem_array[31596] = 16'hbefc;
mem_array[31599] = 16'hea1d;
mem_array[31598] = 16'hbe5e;
mem_array[31601] = 16'h6bb7;
mem_array[31600] = 16'hbe40;
mem_array[31603] = 16'h8bc2;
mem_array[31602] = 16'h3e73;
mem_array[31605] = 16'h0703;
mem_array[31604] = 16'hbf50;
mem_array[31607] = 16'h2abb;
mem_array[31606] = 16'h3d46;
mem_array[31609] = 16'h4dec;
mem_array[31608] = 16'h3b1e;
mem_array[31611] = 16'h0f04;
mem_array[31610] = 16'hbf80;
mem_array[31613] = 16'h02cc;
mem_array[31612] = 16'h3e5e;
mem_array[31615] = 16'h5dc4;
mem_array[31614] = 16'hbe6e;
mem_array[31617] = 16'h12f0;
mem_array[31616] = 16'h3e15;
mem_array[31619] = 16'h715d;
mem_array[31618] = 16'h3e8d;
mem_array[31621] = 16'hcd62;
mem_array[31620] = 16'hbd9d;
mem_array[31623] = 16'h09a8;
mem_array[31622] = 16'hbf2b;
mem_array[31625] = 16'hd8f0;
mem_array[31624] = 16'h3da3;
mem_array[31627] = 16'h7b11;
mem_array[31626] = 16'h3dee;
mem_array[31629] = 16'h0798;
mem_array[31628] = 16'hbe7f;
mem_array[31631] = 16'hb50b;
mem_array[31630] = 16'h3f11;
mem_array[31633] = 16'h7065;
mem_array[31632] = 16'h3d3b;
mem_array[31635] = 16'h51ee;
mem_array[31634] = 16'hbf37;
mem_array[31637] = 16'ha8da;
mem_array[31636] = 16'h3e04;
mem_array[31639] = 16'h90d1;
mem_array[31638] = 16'h3eb6;
mem_array[31641] = 16'hedae;
mem_array[31640] = 16'h3ddd;
mem_array[31643] = 16'hc383;
mem_array[31642] = 16'h3dbb;
mem_array[31645] = 16'hc497;
mem_array[31644] = 16'h3f16;
mem_array[31647] = 16'h2085;
mem_array[31646] = 16'hbd73;
mem_array[31649] = 16'h3da4;
mem_array[31648] = 16'h3d5d;
mem_array[31651] = 16'h33b1;
mem_array[31650] = 16'hbe16;
mem_array[31653] = 16'had02;
mem_array[31652] = 16'h3f03;
mem_array[31655] = 16'hdd96;
mem_array[31654] = 16'h3e5c;
mem_array[31657] = 16'h0952;
mem_array[31656] = 16'hbf76;
mem_array[31659] = 16'h4d87;
mem_array[31658] = 16'h3e08;
mem_array[31661] = 16'h25f4;
mem_array[31660] = 16'h3e94;
mem_array[31663] = 16'h18ea;
mem_array[31662] = 16'h3e91;
mem_array[31665] = 16'hf321;
mem_array[31664] = 16'hbf67;
mem_array[31667] = 16'hffcf;
mem_array[31666] = 16'h3e8b;
mem_array[31669] = 16'h0b3c;
mem_array[31668] = 16'hbf0c;
mem_array[31671] = 16'h8d45;
mem_array[31670] = 16'hbf18;
mem_array[31673] = 16'h05d3;
mem_array[31672] = 16'h3ddd;
mem_array[31675] = 16'h95fb;
mem_array[31674] = 16'hbf35;
mem_array[31677] = 16'hff6f;
mem_array[31676] = 16'h3e54;
mem_array[31679] = 16'hd191;
mem_array[31678] = 16'h3ec2;
mem_array[31681] = 16'h5fc1;
mem_array[31680] = 16'h3e64;
mem_array[31683] = 16'h0dc1;
mem_array[31682] = 16'hbef5;
mem_array[31685] = 16'h3fb6;
mem_array[31684] = 16'h3ee3;
mem_array[31687] = 16'h36cf;
mem_array[31686] = 16'hbdc3;
mem_array[31689] = 16'he829;
mem_array[31688] = 16'hbeda;
mem_array[31691] = 16'h3200;
mem_array[31690] = 16'hbdcf;
mem_array[31693] = 16'h9c0f;
mem_array[31692] = 16'h3c87;
mem_array[31695] = 16'h9988;
mem_array[31694] = 16'h3f1e;
mem_array[31697] = 16'hc85a;
mem_array[31696] = 16'h3ede;
mem_array[31699] = 16'h2c68;
mem_array[31698] = 16'hbe27;
mem_array[31701] = 16'h0a46;
mem_array[31700] = 16'hbd45;
mem_array[31703] = 16'hd3bd;
mem_array[31702] = 16'h3d98;
mem_array[31705] = 16'h67ed;
mem_array[31704] = 16'h3e6e;
mem_array[31707] = 16'hba9c;
mem_array[31706] = 16'hbc99;
mem_array[31709] = 16'heb76;
mem_array[31708] = 16'h3e2f;
mem_array[31711] = 16'h4eaa;
mem_array[31710] = 16'hbe78;
mem_array[31713] = 16'h14b2;
mem_array[31712] = 16'h3e3c;
mem_array[31715] = 16'h5aa6;
mem_array[31714] = 16'h3dee;
mem_array[31717] = 16'ha8c2;
mem_array[31716] = 16'hbfa4;
mem_array[31719] = 16'hcde5;
mem_array[31718] = 16'hbde4;
mem_array[31721] = 16'h4f1f;
mem_array[31720] = 16'h3e93;
mem_array[31723] = 16'h2954;
mem_array[31722] = 16'h3ee7;
mem_array[31725] = 16'h03ff;
mem_array[31724] = 16'hbfb5;
mem_array[31727] = 16'h7763;
mem_array[31726] = 16'h3e6d;
mem_array[31729] = 16'h7315;
mem_array[31728] = 16'h3e23;
mem_array[31731] = 16'h686f;
mem_array[31730] = 16'hbf16;
mem_array[31733] = 16'h5cae;
mem_array[31732] = 16'h3e8f;
mem_array[31735] = 16'h321c;
mem_array[31734] = 16'hbead;
mem_array[31737] = 16'habdd;
mem_array[31736] = 16'h3f00;
mem_array[31739] = 16'hf582;
mem_array[31738] = 16'h3f23;
mem_array[31741] = 16'h8e05;
mem_array[31740] = 16'h3f2c;
mem_array[31743] = 16'h8b53;
mem_array[31742] = 16'h3c24;
mem_array[31745] = 16'hae53;
mem_array[31744] = 16'h3fa1;
mem_array[31747] = 16'h4913;
mem_array[31746] = 16'hbf3a;
mem_array[31749] = 16'h390d;
mem_array[31748] = 16'h3eb6;
mem_array[31751] = 16'h3319;
mem_array[31750] = 16'h3f22;
mem_array[31753] = 16'h72e6;
mem_array[31752] = 16'h3efa;
mem_array[31755] = 16'h7752;
mem_array[31754] = 16'h3f39;
mem_array[31757] = 16'h7789;
mem_array[31756] = 16'h3f85;
mem_array[31759] = 16'h4428;
mem_array[31758] = 16'h3f33;
mem_array[31761] = 16'h1409;
mem_array[31760] = 16'hbd10;
mem_array[31763] = 16'h95ee;
mem_array[31762] = 16'h3cd5;
mem_array[31765] = 16'h20b8;
mem_array[31764] = 16'h3ee8;
mem_array[31767] = 16'h215f;
mem_array[31766] = 16'h3f6f;
mem_array[31769] = 16'h1d16;
mem_array[31768] = 16'h3fa2;
mem_array[31771] = 16'h53bc;
mem_array[31770] = 16'hbdeb;
mem_array[31773] = 16'h358a;
mem_array[31772] = 16'h3f55;
mem_array[31775] = 16'hc8d3;
mem_array[31774] = 16'h3e59;
mem_array[31777] = 16'hd988;
mem_array[31776] = 16'h3dbd;
mem_array[31779] = 16'hd18c;
mem_array[31778] = 16'h3e4c;
mem_array[31781] = 16'hd075;
mem_array[31780] = 16'h3f03;
mem_array[31783] = 16'h73d3;
mem_array[31782] = 16'hbfa5;
mem_array[31785] = 16'h92c0;
mem_array[31784] = 16'hbfbf;
mem_array[31787] = 16'h4d6b;
mem_array[31786] = 16'hbf56;
mem_array[31789] = 16'hf981;
mem_array[31788] = 16'h3f93;
mem_array[31791] = 16'he01b;
mem_array[31790] = 16'h3e90;
mem_array[31793] = 16'h9d3b;
mem_array[31792] = 16'hbf02;
mem_array[31795] = 16'he7de;
mem_array[31794] = 16'hbf03;
mem_array[31797] = 16'h46a7;
mem_array[31796] = 16'h3f2f;
mem_array[31799] = 16'h3cca;
mem_array[31798] = 16'h3df6;
mem_array[31801] = 16'h4be5;
mem_array[31800] = 16'h3f12;
mem_array[31803] = 16'hdb96;
mem_array[31802] = 16'hb9f8;
mem_array[31805] = 16'h60b3;
mem_array[31804] = 16'h3f75;
mem_array[31807] = 16'hdb03;
mem_array[31806] = 16'hbf7b;
mem_array[31809] = 16'hf935;
mem_array[31808] = 16'h3f68;
mem_array[31811] = 16'h5346;
mem_array[31810] = 16'hbd89;
mem_array[31813] = 16'h842c;
mem_array[31812] = 16'h3e8a;
mem_array[31815] = 16'h4c34;
mem_array[31814] = 16'h3e13;
mem_array[31817] = 16'hebf2;
mem_array[31816] = 16'h3f3e;
mem_array[31819] = 16'h97e8;
mem_array[31818] = 16'hbda9;
mem_array[31821] = 16'hadcc;
mem_array[31820] = 16'hbdb2;
mem_array[31823] = 16'ha816;
mem_array[31822] = 16'h3e24;
mem_array[31825] = 16'h7517;
mem_array[31824] = 16'hbf9e;
mem_array[31827] = 16'h850f;
mem_array[31826] = 16'h3f82;
mem_array[31829] = 16'hfd7e;
mem_array[31828] = 16'h3ebc;
mem_array[31831] = 16'hcbdd;
mem_array[31830] = 16'h3e95;
mem_array[31833] = 16'heabc;
mem_array[31832] = 16'h3fa8;
mem_array[31835] = 16'h9409;
mem_array[31834] = 16'hbcc2;
mem_array[31837] = 16'h776c;
mem_array[31836] = 16'h3df0;
mem_array[31839] = 16'h3d12;
mem_array[31838] = 16'h3f1c;
mem_array[31841] = 16'he114;
mem_array[31840] = 16'h3f97;
mem_array[31843] = 16'h2596;
mem_array[31842] = 16'hbe2a;
mem_array[31845] = 16'h4494;
mem_array[31844] = 16'hbea1;
mem_array[31847] = 16'hd72c;
mem_array[31846] = 16'hbf1a;
mem_array[31849] = 16'h1a81;
mem_array[31848] = 16'h3f7c;
mem_array[31851] = 16'hbf93;
mem_array[31850] = 16'h3e61;
mem_array[31853] = 16'hf2a0;
mem_array[31852] = 16'hbd7e;
mem_array[31855] = 16'h1a29;
mem_array[31854] = 16'hbe01;
mem_array[31857] = 16'h5b33;
mem_array[31856] = 16'h3f0a;
mem_array[31859] = 16'haeab;
mem_array[31858] = 16'hbed7;
mem_array[31861] = 16'hbce6;
mem_array[31860] = 16'h3f5e;
mem_array[31863] = 16'h5319;
mem_array[31862] = 16'h3dd5;
mem_array[31865] = 16'hbcf6;
mem_array[31864] = 16'h3e1c;
mem_array[31867] = 16'h7c3b;
mem_array[31866] = 16'hbf19;
mem_array[31869] = 16'h430a;
mem_array[31868] = 16'hbd60;
mem_array[31871] = 16'hebd5;
mem_array[31870] = 16'h3edc;
mem_array[31873] = 16'h454b;
mem_array[31872] = 16'h3f7c;
mem_array[31875] = 16'h2274;
mem_array[31874] = 16'hbe33;
mem_array[31877] = 16'h37c1;
mem_array[31876] = 16'h3f0a;
mem_array[31879] = 16'h0c03;
mem_array[31878] = 16'h3fa9;
mem_array[31881] = 16'hd567;
mem_array[31880] = 16'hbd3f;
mem_array[31883] = 16'h6f01;
mem_array[31882] = 16'hbd6a;
mem_array[31885] = 16'h2573;
mem_array[31884] = 16'hbecf;
mem_array[31887] = 16'h10da;
mem_array[31886] = 16'h3f82;
mem_array[31889] = 16'h1a50;
mem_array[31888] = 16'h3e16;
mem_array[31891] = 16'hea06;
mem_array[31890] = 16'hbf4e;
mem_array[31893] = 16'h01c3;
mem_array[31892] = 16'h3f68;
mem_array[31895] = 16'hb3f6;
mem_array[31894] = 16'h3d7a;
mem_array[31897] = 16'ha7ce;
mem_array[31896] = 16'hbe97;
mem_array[31899] = 16'h750e;
mem_array[31898] = 16'hbe6e;
mem_array[31901] = 16'h0816;
mem_array[31900] = 16'hbee9;
mem_array[31903] = 16'heccc;
mem_array[31902] = 16'hbf05;
mem_array[31905] = 16'hdd99;
mem_array[31904] = 16'hbef3;
mem_array[31907] = 16'h4f77;
mem_array[31906] = 16'hbfa2;
mem_array[31909] = 16'h5f56;
mem_array[31908] = 16'h3e92;
mem_array[31911] = 16'hbdc0;
mem_array[31910] = 16'hbdfb;
mem_array[31913] = 16'h1ffd;
mem_array[31912] = 16'h3f20;
mem_array[31915] = 16'hbca5;
mem_array[31914] = 16'hbe3e;
mem_array[31917] = 16'h7107;
mem_array[31916] = 16'h3eaa;
mem_array[31919] = 16'h296a;
mem_array[31918] = 16'hbf17;
mem_array[31921] = 16'hf272;
mem_array[31920] = 16'h3cf1;
mem_array[31923] = 16'he232;
mem_array[31922] = 16'h3b6a;
mem_array[31925] = 16'hcc01;
mem_array[31924] = 16'hbd3d;
mem_array[31927] = 16'h0373;
mem_array[31926] = 16'h3d6b;
mem_array[31929] = 16'h3c4a;
mem_array[31928] = 16'hbda0;
mem_array[31931] = 16'he69c;
mem_array[31930] = 16'hbcb7;
mem_array[31933] = 16'hf582;
mem_array[31932] = 16'h3cd3;
mem_array[31935] = 16'h6783;
mem_array[31934] = 16'hbd65;
mem_array[31937] = 16'h14bc;
mem_array[31936] = 16'h3c78;
mem_array[31939] = 16'hb661;
mem_array[31938] = 16'h3d88;
mem_array[31941] = 16'h13f2;
mem_array[31940] = 16'hbb82;
mem_array[31943] = 16'h0631;
mem_array[31942] = 16'hbddd;
mem_array[31945] = 16'h02f2;
mem_array[31944] = 16'h3d5a;
mem_array[31947] = 16'h96e7;
mem_array[31946] = 16'hbc34;
mem_array[31949] = 16'h01a4;
mem_array[31948] = 16'h3d05;
mem_array[31951] = 16'hfec3;
mem_array[31950] = 16'h3c94;
mem_array[31953] = 16'hb22b;
mem_array[31952] = 16'h3e24;
mem_array[31955] = 16'h1250;
mem_array[31954] = 16'hbd2e;
mem_array[31957] = 16'hb5e9;
mem_array[31956] = 16'hbd19;
mem_array[31959] = 16'h6700;
mem_array[31958] = 16'hbca1;
mem_array[31961] = 16'hbe4d;
mem_array[31960] = 16'hbdaf;
mem_array[31963] = 16'hcccc;
mem_array[31962] = 16'hbe15;
mem_array[31965] = 16'h36d8;
mem_array[31964] = 16'h3d1b;
mem_array[31967] = 16'h1c35;
mem_array[31966] = 16'hbdfb;
mem_array[31969] = 16'h90db;
mem_array[31968] = 16'hbc72;
mem_array[31971] = 16'hf656;
mem_array[31970] = 16'hbd80;
mem_array[31973] = 16'h7b92;
mem_array[31972] = 16'hbd80;
mem_array[31975] = 16'hd454;
mem_array[31974] = 16'hbde3;
mem_array[31977] = 16'h6303;
mem_array[31976] = 16'hbdb0;
mem_array[31979] = 16'h07dc;
mem_array[31978] = 16'hbca2;
mem_array[31981] = 16'hb53b;
mem_array[31980] = 16'hbd4c;
mem_array[31983] = 16'h699a;
mem_array[31982] = 16'h3f57;
mem_array[31985] = 16'h1ee3;
mem_array[31984] = 16'h3e2c;
mem_array[31987] = 16'hc5c7;
mem_array[31986] = 16'h3d9f;
mem_array[31989] = 16'h8d5a;
mem_array[31988] = 16'hbd10;
mem_array[31991] = 16'h9d7a;
mem_array[31990] = 16'hbdc2;
mem_array[31993] = 16'h49ea;
mem_array[31992] = 16'hbc10;
mem_array[31995] = 16'hd0e4;
mem_array[31994] = 16'hbcba;
mem_array[31997] = 16'h2cf8;
mem_array[31996] = 16'hbc78;
mem_array[31999] = 16'hd28d;
mem_array[31998] = 16'h3e1e;
mem_array[32001] = 16'ha7fb;
mem_array[32000] = 16'hbdbc;
mem_array[32003] = 16'h9cbd;
mem_array[32002] = 16'hbd47;
mem_array[32005] = 16'hec95;
mem_array[32004] = 16'hbd72;
mem_array[32007] = 16'h3cf8;
mem_array[32006] = 16'hbe3f;
mem_array[32009] = 16'hd62d;
mem_array[32008] = 16'h3de8;
mem_array[32011] = 16'hbdb4;
mem_array[32010] = 16'hbf43;
mem_array[32013] = 16'h8984;
mem_array[32012] = 16'hbd22;
mem_array[32015] = 16'h8a49;
mem_array[32014] = 16'hbc42;
mem_array[32017] = 16'h6f55;
mem_array[32016] = 16'hbd69;
mem_array[32019] = 16'h0f25;
mem_array[32018] = 16'h3d4c;
mem_array[32021] = 16'h6fdc;
mem_array[32020] = 16'hbf54;
mem_array[32023] = 16'h0298;
mem_array[32022] = 16'h3f93;
mem_array[32025] = 16'h2777;
mem_array[32024] = 16'h3c08;
mem_array[32027] = 16'h8a83;
mem_array[32026] = 16'hbe23;
mem_array[32029] = 16'hfd41;
mem_array[32028] = 16'hbeff;
mem_array[32031] = 16'h5be5;
mem_array[32030] = 16'h3e8f;
mem_array[32033] = 16'hda29;
mem_array[32032] = 16'h3eab;
mem_array[32035] = 16'heee7;
mem_array[32034] = 16'h3da8;
mem_array[32037] = 16'h18e6;
mem_array[32036] = 16'hbd6b;
mem_array[32039] = 16'h7e72;
mem_array[32038] = 16'hbf71;
mem_array[32041] = 16'h10b9;
mem_array[32040] = 16'h3f00;
mem_array[32043] = 16'he409;
mem_array[32042] = 16'h3f4c;
mem_array[32045] = 16'h9819;
mem_array[32044] = 16'hbdd0;
mem_array[32047] = 16'hbf02;
mem_array[32046] = 16'h3fc6;
mem_array[32049] = 16'h99ac;
mem_array[32048] = 16'hbece;
mem_array[32051] = 16'h5d33;
mem_array[32050] = 16'h3f91;
mem_array[32053] = 16'h7cc0;
mem_array[32052] = 16'hbfaf;
mem_array[32055] = 16'hc757;
mem_array[32054] = 16'hbeea;
mem_array[32057] = 16'h6713;
mem_array[32056] = 16'hbf1c;
mem_array[32059] = 16'h34f3;
mem_array[32058] = 16'hbdd1;
mem_array[32061] = 16'hc051;
mem_array[32060] = 16'hbcec;
mem_array[32063] = 16'h31a5;
mem_array[32062] = 16'hbc8c;
mem_array[32065] = 16'hb50c;
mem_array[32064] = 16'hbdf9;
mem_array[32067] = 16'h5176;
mem_array[32066] = 16'hbef4;
mem_array[32069] = 16'h7edc;
mem_array[32068] = 16'hbf13;
mem_array[32071] = 16'h74a1;
mem_array[32070] = 16'h3e95;
mem_array[32073] = 16'h8f18;
mem_array[32072] = 16'hbf17;
mem_array[32075] = 16'had3c;
mem_array[32074] = 16'hbe8b;
mem_array[32077] = 16'h7200;
mem_array[32076] = 16'h3efd;
mem_array[32079] = 16'h291f;
mem_array[32078] = 16'h3f1a;
mem_array[32081] = 16'h6a0d;
mem_array[32080] = 16'hbf23;
mem_array[32083] = 16'h3395;
mem_array[32082] = 16'h3f1c;
mem_array[32085] = 16'h85c8;
mem_array[32084] = 16'hbe04;
mem_array[32087] = 16'h596f;
mem_array[32086] = 16'hbebd;
mem_array[32089] = 16'h3dfe;
mem_array[32088] = 16'hbeec;
mem_array[32091] = 16'h91a8;
mem_array[32090] = 16'h3f76;
mem_array[32093] = 16'h5dca;
mem_array[32092] = 16'h3fac;
mem_array[32095] = 16'he1b7;
mem_array[32094] = 16'h3ee0;
mem_array[32097] = 16'h1c1e;
mem_array[32096] = 16'h3e8a;
mem_array[32099] = 16'hc9d5;
mem_array[32098] = 16'h3e81;
mem_array[32101] = 16'h1afb;
mem_array[32100] = 16'h3ecc;
mem_array[32103] = 16'hb2cc;
mem_array[32102] = 16'hbf34;
mem_array[32105] = 16'hfb01;
mem_array[32104] = 16'hbf4e;
mem_array[32107] = 16'h1771;
mem_array[32106] = 16'hbeb4;
mem_array[32109] = 16'h3aaa;
mem_array[32108] = 16'h3eec;
mem_array[32111] = 16'had5f;
mem_array[32110] = 16'hbf33;
mem_array[32113] = 16'h4c54;
mem_array[32112] = 16'h3eb3;
mem_array[32115] = 16'h0135;
mem_array[32114] = 16'h3f52;
mem_array[32117] = 16'hb16a;
mem_array[32116] = 16'hbe3c;
mem_array[32119] = 16'h94c6;
mem_array[32118] = 16'hbeb8;
mem_array[32121] = 16'h21ce;
mem_array[32120] = 16'hbb7c;
mem_array[32123] = 16'h038a;
mem_array[32122] = 16'hbbbb;
mem_array[32125] = 16'h07f3;
mem_array[32124] = 16'hbf1b;
mem_array[32127] = 16'h7114;
mem_array[32126] = 16'hbf51;
mem_array[32129] = 16'h5810;
mem_array[32128] = 16'hbdac;
mem_array[32131] = 16'he4f8;
mem_array[32130] = 16'h3e2a;
mem_array[32133] = 16'h6b9b;
mem_array[32132] = 16'h3f27;
mem_array[32135] = 16'h22be;
mem_array[32134] = 16'h3f5e;
mem_array[32137] = 16'h75d1;
mem_array[32136] = 16'hbfd2;
mem_array[32139] = 16'h34ab;
mem_array[32138] = 16'h3ec1;
mem_array[32141] = 16'hc458;
mem_array[32140] = 16'h3f5f;
mem_array[32143] = 16'hbf87;
mem_array[32142] = 16'h3ebb;
mem_array[32145] = 16'h81ea;
mem_array[32144] = 16'hbed4;
mem_array[32147] = 16'h6746;
mem_array[32146] = 16'hbd90;
mem_array[32149] = 16'h7d52;
mem_array[32148] = 16'h3f05;
mem_array[32151] = 16'h59f6;
mem_array[32150] = 16'hbedc;
mem_array[32153] = 16'hf144;
mem_array[32152] = 16'h3e3e;
mem_array[32155] = 16'hd10f;
mem_array[32154] = 16'h3e16;
mem_array[32157] = 16'h04bd;
mem_array[32156] = 16'h3d71;
mem_array[32159] = 16'h8c99;
mem_array[32158] = 16'h3f4e;
mem_array[32161] = 16'h997f;
mem_array[32160] = 16'h3d25;
mem_array[32163] = 16'h716c;
mem_array[32162] = 16'hbd8a;
mem_array[32165] = 16'h3c0e;
mem_array[32164] = 16'hbdc1;
mem_array[32167] = 16'h8712;
mem_array[32166] = 16'hbd29;
mem_array[32169] = 16'haada;
mem_array[32168] = 16'h3da6;
mem_array[32171] = 16'h14b2;
mem_array[32170] = 16'hbe74;
mem_array[32173] = 16'h86e1;
mem_array[32172] = 16'hbe84;
mem_array[32175] = 16'h7778;
mem_array[32174] = 16'h3c8c;
mem_array[32177] = 16'h26db;
mem_array[32176] = 16'h3ec8;
mem_array[32179] = 16'hc70a;
mem_array[32178] = 16'hbdac;
mem_array[32181] = 16'h654e;
mem_array[32180] = 16'h3d3e;
mem_array[32183] = 16'h52cf;
mem_array[32182] = 16'h3da1;
mem_array[32185] = 16'h5745;
mem_array[32184] = 16'h3e7e;
mem_array[32187] = 16'h3c63;
mem_array[32186] = 16'hbe41;
mem_array[32189] = 16'h01c1;
mem_array[32188] = 16'hbe08;
mem_array[32191] = 16'he848;
mem_array[32190] = 16'hbd8c;
mem_array[32193] = 16'h7aed;
mem_array[32192] = 16'h3f3a;
mem_array[32195] = 16'hf679;
mem_array[32194] = 16'h3d77;
mem_array[32197] = 16'h2f18;
mem_array[32196] = 16'hbffc;
mem_array[32199] = 16'h77f2;
mem_array[32198] = 16'hbdac;
mem_array[32201] = 16'hbf1b;
mem_array[32200] = 16'h3f5e;
mem_array[32203] = 16'h5b9c;
mem_array[32202] = 16'hbd42;
mem_array[32205] = 16'he3c2;
mem_array[32204] = 16'hbf58;
mem_array[32207] = 16'h9553;
mem_array[32206] = 16'h3e43;
mem_array[32209] = 16'hb376;
mem_array[32208] = 16'h3e75;
mem_array[32211] = 16'h5b0e;
mem_array[32210] = 16'hbe8b;
mem_array[32213] = 16'hc8a2;
mem_array[32212] = 16'h3e0b;
mem_array[32215] = 16'h3196;
mem_array[32214] = 16'h3f08;
mem_array[32217] = 16'hbc57;
mem_array[32216] = 16'hbd88;
mem_array[32219] = 16'h7c23;
mem_array[32218] = 16'h3e0d;
mem_array[32221] = 16'hb3e8;
mem_array[32220] = 16'hbf81;
mem_array[32223] = 16'hec26;
mem_array[32222] = 16'hbe52;
mem_array[32225] = 16'h59c1;
mem_array[32224] = 16'hbeb8;
mem_array[32227] = 16'hfdb2;
mem_array[32226] = 16'h3ebc;
mem_array[32229] = 16'h3309;
mem_array[32228] = 16'h3db2;
mem_array[32231] = 16'h25c0;
mem_array[32230] = 16'h3e22;
mem_array[32233] = 16'h712b;
mem_array[32232] = 16'h3ead;
mem_array[32235] = 16'h03a1;
mem_array[32234] = 16'hbdb3;
mem_array[32237] = 16'h85b6;
mem_array[32236] = 16'h3eb7;
mem_array[32239] = 16'hefcf;
mem_array[32238] = 16'hbe4d;
mem_array[32241] = 16'h4401;
mem_array[32240] = 16'hbd8a;
mem_array[32243] = 16'h0ae2;
mem_array[32242] = 16'hbdb3;
mem_array[32245] = 16'hab5a;
mem_array[32244] = 16'hbccb;
mem_array[32247] = 16'he244;
mem_array[32246] = 16'h3d2a;
mem_array[32249] = 16'h63b7;
mem_array[32248] = 16'hbdcd;
mem_array[32251] = 16'hd400;
mem_array[32250] = 16'hbe9d;
mem_array[32253] = 16'h4387;
mem_array[32252] = 16'h3df4;
mem_array[32255] = 16'h792e;
mem_array[32254] = 16'hbcd5;
mem_array[32257] = 16'h2efc;
mem_array[32256] = 16'hbf38;
mem_array[32259] = 16'h6de0;
mem_array[32258] = 16'h3e18;
mem_array[32261] = 16'h5c10;
mem_array[32260] = 16'hbe4e;
mem_array[32263] = 16'hc5b5;
mem_array[32262] = 16'hbdc9;
mem_array[32265] = 16'h68d6;
mem_array[32264] = 16'hbfa6;
mem_array[32267] = 16'h7eeb;
mem_array[32266] = 16'h3c8d;
mem_array[32269] = 16'he900;
mem_array[32268] = 16'h3e95;
mem_array[32271] = 16'hfc01;
mem_array[32270] = 16'hbcab;
mem_array[32273] = 16'hd192;
mem_array[32272] = 16'h3ca6;
mem_array[32275] = 16'h56e0;
mem_array[32274] = 16'h3eda;
mem_array[32277] = 16'hc5d2;
mem_array[32276] = 16'h3e68;
mem_array[32279] = 16'ha3ab;
mem_array[32278] = 16'hbed6;
mem_array[32281] = 16'hf1b7;
mem_array[32280] = 16'hbf05;
mem_array[32283] = 16'hcec5;
mem_array[32282] = 16'hbe67;
mem_array[32285] = 16'h8e80;
mem_array[32284] = 16'hbdb8;
mem_array[32287] = 16'h10a1;
mem_array[32286] = 16'h3e15;
mem_array[32289] = 16'h10cf;
mem_array[32288] = 16'hbeff;
mem_array[32291] = 16'hd096;
mem_array[32290] = 16'h3e37;
mem_array[32293] = 16'h90a0;
mem_array[32292] = 16'hbb24;
mem_array[32295] = 16'h60a8;
mem_array[32294] = 16'hbe08;
mem_array[32297] = 16'h8ce7;
mem_array[32296] = 16'hbd3f;
mem_array[32299] = 16'ha71e;
mem_array[32298] = 16'hbfa4;
mem_array[32301] = 16'h610c;
mem_array[32300] = 16'h3c43;
mem_array[32303] = 16'h0b5a;
mem_array[32302] = 16'h3d1c;
mem_array[32305] = 16'hd8d7;
mem_array[32304] = 16'hbcba;
mem_array[32307] = 16'he298;
mem_array[32306] = 16'h3d6c;
mem_array[32309] = 16'h1418;
mem_array[32308] = 16'h3ec6;
mem_array[32311] = 16'hb22a;
mem_array[32310] = 16'h3d20;
mem_array[32313] = 16'hfe4b;
mem_array[32312] = 16'hbee4;
mem_array[32315] = 16'hf787;
mem_array[32314] = 16'h3e28;
mem_array[32317] = 16'h07ce;
mem_array[32316] = 16'hbe2d;
mem_array[32319] = 16'heb96;
mem_array[32318] = 16'h3ecd;
mem_array[32321] = 16'h4ed1;
mem_array[32320] = 16'hbedf;
mem_array[32323] = 16'ha9d8;
mem_array[32322] = 16'h3e9f;
mem_array[32325] = 16'hec01;
mem_array[32324] = 16'h3dcc;
mem_array[32327] = 16'h7482;
mem_array[32326] = 16'h3e15;
mem_array[32329] = 16'h7b7a;
mem_array[32328] = 16'hbde5;
mem_array[32331] = 16'h8a2b;
mem_array[32330] = 16'hbf2f;
mem_array[32333] = 16'h56e2;
mem_array[32332] = 16'h3e32;
mem_array[32335] = 16'h58cc;
mem_array[32334] = 16'h3ed5;
mem_array[32337] = 16'heb08;
mem_array[32336] = 16'hbdf6;
mem_array[32339] = 16'hf8fb;
mem_array[32338] = 16'hbea6;
mem_array[32341] = 16'h3348;
mem_array[32340] = 16'h3e4a;
mem_array[32343] = 16'h40df;
mem_array[32342] = 16'hbd3b;
mem_array[32345] = 16'h1921;
mem_array[32344] = 16'h3e6e;
mem_array[32347] = 16'hedcc;
mem_array[32346] = 16'h3e85;
mem_array[32349] = 16'h4753;
mem_array[32348] = 16'hbe96;
mem_array[32351] = 16'h248f;
mem_array[32350] = 16'h3daa;
mem_array[32353] = 16'hc535;
mem_array[32352] = 16'h3e84;
mem_array[32355] = 16'hd766;
mem_array[32354] = 16'hbd06;
mem_array[32357] = 16'h3cc9;
mem_array[32356] = 16'h3d92;
mem_array[32359] = 16'h1ffc;
mem_array[32358] = 16'hbea2;
mem_array[32361] = 16'h2544;
mem_array[32360] = 16'hbc9a;
mem_array[32363] = 16'h45fb;
mem_array[32362] = 16'hbd5f;
mem_array[32365] = 16'h8058;
mem_array[32364] = 16'h3e06;
mem_array[32367] = 16'ha877;
mem_array[32366] = 16'h3e73;
mem_array[32369] = 16'hc024;
mem_array[32368] = 16'h3f1c;
mem_array[32371] = 16'h6fb5;
mem_array[32370] = 16'h3e64;
mem_array[32373] = 16'hdbc5;
mem_array[32372] = 16'hbdcd;
mem_array[32375] = 16'h48e2;
mem_array[32374] = 16'hbea0;
mem_array[32377] = 16'h98fe;
mem_array[32376] = 16'h3eb4;
mem_array[32379] = 16'h2074;
mem_array[32378] = 16'h3e50;
mem_array[32381] = 16'h1927;
mem_array[32380] = 16'hbfbf;
mem_array[32383] = 16'h33b4;
mem_array[32382] = 16'h3dcd;
mem_array[32385] = 16'h5f91;
mem_array[32384] = 16'h3e17;
mem_array[32387] = 16'hb53d;
mem_array[32386] = 16'h3e45;
mem_array[32389] = 16'h4d58;
mem_array[32388] = 16'hbebe;
mem_array[32391] = 16'h07da;
mem_array[32390] = 16'h3e0b;
mem_array[32393] = 16'hd74f;
mem_array[32392] = 16'hbcec;
mem_array[32395] = 16'h352d;
mem_array[32394] = 16'h3e5f;
mem_array[32397] = 16'h930c;
mem_array[32396] = 16'hbd73;
mem_array[32399] = 16'h59e2;
mem_array[32398] = 16'h3c80;
mem_array[32401] = 16'h1c97;
mem_array[32400] = 16'h3da7;
mem_array[32403] = 16'hbf47;
mem_array[32402] = 16'hbf07;
mem_array[32405] = 16'h8f21;
mem_array[32404] = 16'h3c7a;
mem_array[32407] = 16'hdd57;
mem_array[32406] = 16'h3e8b;
mem_array[32409] = 16'hd51a;
mem_array[32408] = 16'hbec0;
mem_array[32411] = 16'h5593;
mem_array[32410] = 16'h3e7b;
mem_array[32413] = 16'h669d;
mem_array[32412] = 16'h3e5d;
mem_array[32415] = 16'h85d3;
mem_array[32414] = 16'h3dd9;
mem_array[32417] = 16'h9cca;
mem_array[32416] = 16'hbd8b;
mem_array[32419] = 16'h9402;
mem_array[32418] = 16'hbf06;
mem_array[32421] = 16'h4332;
mem_array[32420] = 16'h3c65;
mem_array[32423] = 16'h36e2;
mem_array[32422] = 16'hbcae;
mem_array[32425] = 16'h7d68;
mem_array[32424] = 16'h3e88;
mem_array[32427] = 16'he743;
mem_array[32426] = 16'h3e1b;
mem_array[32429] = 16'hf997;
mem_array[32428] = 16'h3e71;
mem_array[32431] = 16'h7cd6;
mem_array[32430] = 16'h3e7c;
mem_array[32433] = 16'h8566;
mem_array[32432] = 16'hbd49;
mem_array[32435] = 16'h8b32;
mem_array[32434] = 16'hbdc7;
mem_array[32437] = 16'hfab4;
mem_array[32436] = 16'hbd67;
mem_array[32439] = 16'h36e5;
mem_array[32438] = 16'h3ed5;
mem_array[32441] = 16'h0a36;
mem_array[32440] = 16'hbfcc;
mem_array[32443] = 16'h6d48;
mem_array[32442] = 16'h3ea0;
mem_array[32445] = 16'hcaae;
mem_array[32444] = 16'h3da0;
mem_array[32447] = 16'h3128;
mem_array[32446] = 16'h3f0e;
mem_array[32449] = 16'hf7ab;
mem_array[32448] = 16'hbeda;
mem_array[32451] = 16'hb9f1;
mem_array[32450] = 16'hbdc5;
mem_array[32453] = 16'h99c5;
mem_array[32452] = 16'hbd3c;
mem_array[32455] = 16'hb138;
mem_array[32454] = 16'h3d20;
mem_array[32457] = 16'hbd76;
mem_array[32456] = 16'hbe07;
mem_array[32459] = 16'h47da;
mem_array[32458] = 16'h3e30;
mem_array[32461] = 16'h0398;
mem_array[32460] = 16'h3e11;
mem_array[32463] = 16'h9d92;
mem_array[32462] = 16'hbf98;
mem_array[32465] = 16'h2dd5;
mem_array[32464] = 16'hbc8f;
mem_array[32467] = 16'h5a19;
mem_array[32466] = 16'h3f53;
mem_array[32469] = 16'h241a;
mem_array[32468] = 16'hbe08;
mem_array[32471] = 16'h83bc;
mem_array[32470] = 16'h3eb4;
mem_array[32473] = 16'h2700;
mem_array[32472] = 16'h3e16;
mem_array[32475] = 16'h7e13;
mem_array[32474] = 16'h3e99;
mem_array[32477] = 16'h4d6a;
mem_array[32476] = 16'h3ca6;
mem_array[32479] = 16'h2a66;
mem_array[32478] = 16'h3e92;
mem_array[32481] = 16'h5d15;
mem_array[32480] = 16'hbc7c;
mem_array[32483] = 16'hb46f;
mem_array[32482] = 16'hbd4d;
mem_array[32485] = 16'he6de;
mem_array[32484] = 16'h3e9a;
mem_array[32487] = 16'h4b0f;
mem_array[32486] = 16'h3e26;
mem_array[32489] = 16'h080d;
mem_array[32488] = 16'h3e62;
mem_array[32491] = 16'hdd17;
mem_array[32490] = 16'h3ec8;
mem_array[32493] = 16'he9e3;
mem_array[32492] = 16'h3e7e;
mem_array[32495] = 16'hf652;
mem_array[32494] = 16'hbe6d;
mem_array[32497] = 16'h59b1;
mem_array[32496] = 16'hbd3e;
mem_array[32499] = 16'h05b5;
mem_array[32498] = 16'h3e8e;
mem_array[32501] = 16'h1a02;
mem_array[32500] = 16'hbf93;
mem_array[32503] = 16'hc72f;
mem_array[32502] = 16'hbc66;
mem_array[32505] = 16'h9130;
mem_array[32504] = 16'h3ec0;
mem_array[32507] = 16'h94fe;
mem_array[32506] = 16'h3e5c;
mem_array[32509] = 16'h858f;
mem_array[32508] = 16'hbe91;
mem_array[32511] = 16'hddce;
mem_array[32510] = 16'hbc91;
mem_array[32513] = 16'ha906;
mem_array[32512] = 16'hbe4d;
mem_array[32515] = 16'h232e;
mem_array[32514] = 16'hbd32;
mem_array[32517] = 16'h79ca;
mem_array[32516] = 16'hbe0b;
mem_array[32519] = 16'h50a7;
mem_array[32518] = 16'h3ebe;
mem_array[32521] = 16'h3149;
mem_array[32520] = 16'h3ece;
mem_array[32523] = 16'h3574;
mem_array[32522] = 16'hbfa8;
mem_array[32525] = 16'haa86;
mem_array[32524] = 16'h3d41;
mem_array[32527] = 16'hda50;
mem_array[32526] = 16'h3f0a;
mem_array[32529] = 16'ha474;
mem_array[32528] = 16'hbdf2;
mem_array[32531] = 16'h5ae7;
mem_array[32530] = 16'h3ea8;
mem_array[32533] = 16'h5df7;
mem_array[32532] = 16'h3f0b;
mem_array[32535] = 16'h0837;
mem_array[32534] = 16'h3e3b;
mem_array[32537] = 16'h89a0;
mem_array[32536] = 16'h3eac;
mem_array[32539] = 16'h7956;
mem_array[32538] = 16'hbe11;
mem_array[32541] = 16'hffe0;
mem_array[32540] = 16'hbd50;
mem_array[32543] = 16'h30dc;
mem_array[32542] = 16'h3d36;
mem_array[32545] = 16'hdf0a;
mem_array[32544] = 16'h3f28;
mem_array[32547] = 16'h4c41;
mem_array[32546] = 16'h3ddf;
mem_array[32549] = 16'h8a34;
mem_array[32548] = 16'h3ce1;
mem_array[32551] = 16'h22d0;
mem_array[32550] = 16'h3f23;
mem_array[32553] = 16'h7482;
mem_array[32552] = 16'h3eda;
mem_array[32555] = 16'h4afa;
mem_array[32554] = 16'hbe5d;
mem_array[32557] = 16'h9701;
mem_array[32556] = 16'hbe70;
mem_array[32559] = 16'hce75;
mem_array[32558] = 16'hbdbf;
mem_array[32561] = 16'hcc16;
mem_array[32560] = 16'hbf37;
mem_array[32563] = 16'h89ce;
mem_array[32562] = 16'h3e53;
mem_array[32565] = 16'h2f87;
mem_array[32564] = 16'h3eec;
mem_array[32567] = 16'h9734;
mem_array[32566] = 16'h3f16;
mem_array[32569] = 16'h1ae3;
mem_array[32568] = 16'hbf08;
mem_array[32571] = 16'h2bcd;
mem_array[32570] = 16'hbe47;
mem_array[32573] = 16'h615d;
mem_array[32572] = 16'hbd51;
mem_array[32575] = 16'h27a1;
mem_array[32574] = 16'hbc26;
mem_array[32577] = 16'h602b;
mem_array[32576] = 16'hbceb;
mem_array[32579] = 16'he5e5;
mem_array[32578] = 16'h3ea8;
mem_array[32581] = 16'ha356;
mem_array[32580] = 16'h3f05;
mem_array[32583] = 16'h9811;
mem_array[32582] = 16'hbdca;
mem_array[32585] = 16'hb801;
mem_array[32584] = 16'h3e9e;
mem_array[32587] = 16'h938c;
mem_array[32586] = 16'h3d3a;
mem_array[32589] = 16'h6b2f;
mem_array[32588] = 16'h3e6b;
mem_array[32591] = 16'h7f24;
mem_array[32590] = 16'h3e94;
mem_array[32593] = 16'h2691;
mem_array[32592] = 16'h3f28;
mem_array[32595] = 16'h9a37;
mem_array[32594] = 16'h3e84;
mem_array[32597] = 16'hb4f7;
mem_array[32596] = 16'h3d81;
mem_array[32599] = 16'ha328;
mem_array[32598] = 16'hbe70;
mem_array[32601] = 16'h6c75;
mem_array[32600] = 16'hbcdb;
mem_array[32603] = 16'hcbaa;
mem_array[32602] = 16'h3cec;
mem_array[32605] = 16'ha02a;
mem_array[32604] = 16'h3ee3;
mem_array[32607] = 16'hfa9f;
mem_array[32606] = 16'h3df9;
mem_array[32609] = 16'hf821;
mem_array[32608] = 16'h3dff;
mem_array[32611] = 16'h4d2c;
mem_array[32610] = 16'h3f28;
mem_array[32613] = 16'hdaf4;
mem_array[32612] = 16'h3ef1;
mem_array[32615] = 16'hfccf;
mem_array[32614] = 16'hbe38;
mem_array[32617] = 16'h2188;
mem_array[32616] = 16'h3b75;
mem_array[32619] = 16'hf076;
mem_array[32618] = 16'hbe64;
mem_array[32621] = 16'hfe63;
mem_array[32620] = 16'hbdb6;
mem_array[32623] = 16'h7f37;
mem_array[32622] = 16'h3ea0;
mem_array[32625] = 16'hf8e7;
mem_array[32624] = 16'h3f2f;
mem_array[32627] = 16'h5593;
mem_array[32626] = 16'h3f35;
mem_array[32629] = 16'h574f;
mem_array[32628] = 16'hbe8d;
mem_array[32631] = 16'h26fc;
mem_array[32630] = 16'hbe45;
mem_array[32633] = 16'h92e1;
mem_array[32632] = 16'hbcbd;
mem_array[32635] = 16'hdabd;
mem_array[32634] = 16'hbc8f;
mem_array[32637] = 16'h2214;
mem_array[32636] = 16'hbe50;
mem_array[32639] = 16'h6f55;
mem_array[32638] = 16'h3e5c;
mem_array[32641] = 16'hda6e;
mem_array[32640] = 16'h3eaf;
mem_array[32643] = 16'ha861;
mem_array[32642] = 16'h3e79;
mem_array[32645] = 16'hfbc5;
mem_array[32644] = 16'h3edb;
mem_array[32647] = 16'h5182;
mem_array[32646] = 16'hbe6d;
mem_array[32649] = 16'h8c94;
mem_array[32648] = 16'h3ec9;
mem_array[32651] = 16'h2bc3;
mem_array[32650] = 16'hbb16;
mem_array[32653] = 16'h7316;
mem_array[32652] = 16'h3edf;
mem_array[32655] = 16'haaa9;
mem_array[32654] = 16'h3efc;
mem_array[32657] = 16'h08c2;
mem_array[32656] = 16'hbe8b;
mem_array[32659] = 16'hc089;
mem_array[32658] = 16'h3d7b;
mem_array[32661] = 16'h0aa1;
mem_array[32660] = 16'hbb27;
mem_array[32663] = 16'h1ebe;
mem_array[32662] = 16'hbd5f;
mem_array[32665] = 16'h28fc;
mem_array[32664] = 16'h3ea4;
mem_array[32667] = 16'hea6a;
mem_array[32666] = 16'hbdc7;
mem_array[32669] = 16'h87c8;
mem_array[32668] = 16'h3e33;
mem_array[32671] = 16'hbbfa;
mem_array[32670] = 16'h3f05;
mem_array[32673] = 16'h58cc;
mem_array[32672] = 16'h3e9b;
mem_array[32675] = 16'hf2cf;
mem_array[32674] = 16'hbed4;
mem_array[32677] = 16'h997e;
mem_array[32676] = 16'h3e1d;
mem_array[32679] = 16'hf5d0;
mem_array[32678] = 16'hbea8;
mem_array[32681] = 16'hb149;
mem_array[32680] = 16'hbeec;
mem_array[32683] = 16'hde09;
mem_array[32682] = 16'h3ecd;
mem_array[32685] = 16'habe8;
mem_array[32684] = 16'h3f40;
mem_array[32687] = 16'hdc63;
mem_array[32686] = 16'h3f28;
mem_array[32689] = 16'hec6c;
mem_array[32688] = 16'hbedb;
mem_array[32691] = 16'h6a58;
mem_array[32690] = 16'hbddd;
mem_array[32693] = 16'h8660;
mem_array[32692] = 16'h3e53;
mem_array[32695] = 16'h0d1f;
mem_array[32694] = 16'h3eb2;
mem_array[32697] = 16'h856d;
mem_array[32696] = 16'hbeb3;
mem_array[32699] = 16'hfe43;
mem_array[32698] = 16'h3e53;
mem_array[32701] = 16'haf49;
mem_array[32700] = 16'h3e1e;
mem_array[32703] = 16'h8f3f;
mem_array[32702] = 16'h3e49;
mem_array[32705] = 16'h1972;
mem_array[32704] = 16'h3f03;
mem_array[32707] = 16'h3e03;
mem_array[32706] = 16'hbe60;
mem_array[32709] = 16'hcfc5;
mem_array[32708] = 16'hbd47;
mem_array[32711] = 16'h7ab1;
mem_array[32710] = 16'h3e0a;
mem_array[32713] = 16'hfb8b;
mem_array[32712] = 16'h3df0;
mem_array[32715] = 16'h1722;
mem_array[32714] = 16'h3e5a;
mem_array[32717] = 16'h7a64;
mem_array[32716] = 16'hbe51;
mem_array[32719] = 16'h9479;
mem_array[32718] = 16'h3eb6;
mem_array[32721] = 16'hd028;
mem_array[32720] = 16'hbe11;
mem_array[32723] = 16'hc47a;
mem_array[32722] = 16'hbcd0;
mem_array[32725] = 16'h4704;
mem_array[32724] = 16'h3ea5;
mem_array[32727] = 16'hc2ca;
mem_array[32726] = 16'hbbd5;
mem_array[32729] = 16'h6892;
mem_array[32728] = 16'h3eb6;
mem_array[32731] = 16'hbc1a;
mem_array[32730] = 16'h3eb4;
mem_array[32733] = 16'hc635;
mem_array[32732] = 16'h3dac;
mem_array[32735] = 16'h2c06;
mem_array[32734] = 16'hbdea;
mem_array[32737] = 16'hd552;
mem_array[32736] = 16'hbe29;
mem_array[32739] = 16'h4c5d;
mem_array[32738] = 16'h3d81;
mem_array[32741] = 16'h7bdb;
mem_array[32740] = 16'hbe9b;
mem_array[32743] = 16'h91ed;
mem_array[32742] = 16'h3e84;
mem_array[32745] = 16'h6b07;
mem_array[32744] = 16'hbcdf;
mem_array[32747] = 16'hfe14;
mem_array[32746] = 16'h3e8e;
mem_array[32749] = 16'h2b2c;
mem_array[32748] = 16'hbe21;
mem_array[32751] = 16'h1669;
mem_array[32750] = 16'hbdee;
mem_array[32753] = 16'h2bc8;
mem_array[32752] = 16'h3e04;
mem_array[32755] = 16'h093c;
mem_array[32754] = 16'h3eda;
mem_array[32757] = 16'h0303;
mem_array[32756] = 16'hbe9a;
mem_array[32759] = 16'h2ced;
mem_array[32758] = 16'h3e66;
mem_array[32761] = 16'hb939;
mem_array[32760] = 16'hbef6;
mem_array[32763] = 16'h03c9;
mem_array[32762] = 16'h3eec;
mem_array[32765] = 16'h3477;
mem_array[32764] = 16'h3e88;
mem_array[32767] = 16'h7ba0;
mem_array[32766] = 16'hbb15;
mem_array[32769] = 16'h05b4;
mem_array[32768] = 16'hbee6;
mem_array[32771] = 16'h7353;
mem_array[32770] = 16'h3eb0;
mem_array[32773] = 16'h86f4;
mem_array[32772] = 16'h3dbc;
mem_array[32775] = 16'h7ca8;
mem_array[32774] = 16'hbd39;
mem_array[32777] = 16'h2fab;
mem_array[32776] = 16'h3d79;
mem_array[32779] = 16'hd934;
mem_array[32778] = 16'h3ee8;
mem_array[32781] = 16'h7c0d;
mem_array[32780] = 16'hbd48;
mem_array[32783] = 16'hab73;
mem_array[32782] = 16'h3b9b;
mem_array[32785] = 16'h2619;
mem_array[32784] = 16'h3ef4;
mem_array[32787] = 16'hdfc6;
mem_array[32786] = 16'h3da4;
mem_array[32789] = 16'h221d;
mem_array[32788] = 16'h3e77;
mem_array[32791] = 16'h7e89;
mem_array[32790] = 16'h3d22;
mem_array[32793] = 16'h2348;
mem_array[32792] = 16'hbeb9;
mem_array[32795] = 16'hd0d5;
mem_array[32794] = 16'hbd0e;
mem_array[32797] = 16'hd355;
mem_array[32796] = 16'h3e87;
mem_array[32799] = 16'h6855;
mem_array[32798] = 16'h3e4e;
mem_array[32801] = 16'h25a4;
mem_array[32800] = 16'hbd42;
mem_array[32803] = 16'h9d88;
mem_array[32802] = 16'hbdb5;
mem_array[32805] = 16'hc13b;
mem_array[32804] = 16'h3cec;
mem_array[32807] = 16'h1cd9;
mem_array[32806] = 16'h3e6a;
mem_array[32809] = 16'hb9c3;
mem_array[32808] = 16'h3e02;
mem_array[32811] = 16'h489b;
mem_array[32810] = 16'h3e25;
mem_array[32813] = 16'h603f;
mem_array[32812] = 16'hbec4;
mem_array[32815] = 16'h3af6;
mem_array[32814] = 16'hbdba;
mem_array[32817] = 16'hf3ca;
mem_array[32816] = 16'hbf0b;
mem_array[32819] = 16'hd754;
mem_array[32818] = 16'h3ded;
mem_array[32821] = 16'h8533;
mem_array[32820] = 16'hbee6;
mem_array[32823] = 16'h311c;
mem_array[32822] = 16'hbdee;
mem_array[32825] = 16'hfd1d;
mem_array[32824] = 16'hbcca;
mem_array[32827] = 16'he305;
mem_array[32826] = 16'hbe02;
mem_array[32829] = 16'hb826;
mem_array[32828] = 16'hbe95;
mem_array[32831] = 16'ha9c4;
mem_array[32830] = 16'h3e03;
mem_array[32833] = 16'hcbdf;
mem_array[32832] = 16'hbe08;
mem_array[32835] = 16'h49d4;
mem_array[32834] = 16'h3d92;
mem_array[32837] = 16'hfa18;
mem_array[32836] = 16'hbdef;
mem_array[32839] = 16'hb07b;
mem_array[32838] = 16'h3dd7;
mem_array[32841] = 16'h59de;
mem_array[32840] = 16'hbd96;
mem_array[32843] = 16'h4325;
mem_array[32842] = 16'hbc25;
mem_array[32845] = 16'hb4c4;
mem_array[32844] = 16'h3e1e;
mem_array[32847] = 16'h614b;
mem_array[32846] = 16'h3eab;
mem_array[32849] = 16'hf524;
mem_array[32848] = 16'h3d4f;
mem_array[32851] = 16'hef10;
mem_array[32850] = 16'hbd8a;
mem_array[32853] = 16'h9065;
mem_array[32852] = 16'hbf2e;
mem_array[32855] = 16'h2c37;
mem_array[32854] = 16'hbd7d;
mem_array[32857] = 16'h382f;
mem_array[32856] = 16'h3e5f;
mem_array[32859] = 16'hd078;
mem_array[32858] = 16'h3e62;
mem_array[32861] = 16'h5530;
mem_array[32860] = 16'hbe1e;
mem_array[32863] = 16'hea24;
mem_array[32862] = 16'h3dc8;
mem_array[32865] = 16'h38db;
mem_array[32864] = 16'h3eb8;
mem_array[32867] = 16'h9e91;
mem_array[32866] = 16'h3c94;
mem_array[32869] = 16'h343c;
mem_array[32868] = 16'hbd1f;
mem_array[32871] = 16'he2ab;
mem_array[32870] = 16'hbe16;
mem_array[32873] = 16'he350;
mem_array[32872] = 16'hbd25;
mem_array[32875] = 16'h5f27;
mem_array[32874] = 16'h3e9d;
mem_array[32877] = 16'hf90d;
mem_array[32876] = 16'hbe74;
mem_array[32879] = 16'h522c;
mem_array[32878] = 16'h3e89;
mem_array[32881] = 16'h3248;
mem_array[32880] = 16'hbf1f;
mem_array[32883] = 16'hd1fc;
mem_array[32882] = 16'hbdb9;
mem_array[32885] = 16'h2ef5;
mem_array[32884] = 16'hbde6;
mem_array[32887] = 16'h753c;
mem_array[32886] = 16'hbd98;
mem_array[32889] = 16'h5d91;
mem_array[32888] = 16'hbe53;
mem_array[32891] = 16'h5cf8;
mem_array[32890] = 16'h3e16;
mem_array[32893] = 16'ha249;
mem_array[32892] = 16'hbdf3;
mem_array[32895] = 16'h8bde;
mem_array[32894] = 16'h3cbb;
mem_array[32897] = 16'h05e8;
mem_array[32896] = 16'h3e0d;
mem_array[32899] = 16'hdcc3;
mem_array[32898] = 16'hbae8;
mem_array[32901] = 16'hd2cf;
mem_array[32900] = 16'hbd26;
mem_array[32903] = 16'hc6a5;
mem_array[32902] = 16'h3cd0;
mem_array[32905] = 16'h3fb0;
mem_array[32904] = 16'h3e14;
mem_array[32907] = 16'h6ebe;
mem_array[32906] = 16'h3e47;
mem_array[32909] = 16'h5466;
mem_array[32908] = 16'hbe02;
mem_array[32911] = 16'h8193;
mem_array[32910] = 16'hbdf5;
mem_array[32913] = 16'h3d56;
mem_array[32912] = 16'hbcf8;
mem_array[32915] = 16'h4d67;
mem_array[32914] = 16'hbcec;
mem_array[32917] = 16'had45;
mem_array[32916] = 16'hbdcc;
mem_array[32919] = 16'hc1ef;
mem_array[32918] = 16'h3e7f;
mem_array[32921] = 16'hf933;
mem_array[32920] = 16'hbe95;
mem_array[32923] = 16'hebf7;
mem_array[32922] = 16'h3e29;
mem_array[32925] = 16'h28ca;
mem_array[32924] = 16'h3e3c;
mem_array[32927] = 16'h65b6;
mem_array[32926] = 16'h3e04;
mem_array[32929] = 16'h8b81;
mem_array[32928] = 16'h3d30;
mem_array[32931] = 16'hd574;
mem_array[32930] = 16'hbedc;
mem_array[32933] = 16'h46ec;
mem_array[32932] = 16'h3d95;
mem_array[32935] = 16'h9136;
mem_array[32934] = 16'h3ed1;
mem_array[32937] = 16'h96fd;
mem_array[32936] = 16'hbdff;
mem_array[32939] = 16'hf660;
mem_array[32938] = 16'h3bcd;
mem_array[32941] = 16'h1c82;
mem_array[32940] = 16'h3eb3;
mem_array[32943] = 16'hfa81;
mem_array[32942] = 16'h3d68;
mem_array[32945] = 16'h319d;
mem_array[32944] = 16'hbe13;
mem_array[32947] = 16'ha0c5;
mem_array[32946] = 16'h3dad;
mem_array[32949] = 16'h5e77;
mem_array[32948] = 16'hbe41;
mem_array[32951] = 16'h51ac;
mem_array[32950] = 16'hbdf2;
mem_array[32953] = 16'h8cf2;
mem_array[32952] = 16'h3e1d;
mem_array[32955] = 16'h1db0;
mem_array[32954] = 16'h3d8e;
mem_array[32957] = 16'hb93a;
mem_array[32956] = 16'h3e39;
mem_array[32959] = 16'hce63;
mem_array[32958] = 16'hbda6;
mem_array[32961] = 16'h0791;
mem_array[32960] = 16'hbd43;
mem_array[32963] = 16'hb7d4;
mem_array[32962] = 16'h3d93;
mem_array[32965] = 16'h6df2;
mem_array[32964] = 16'h3e00;
mem_array[32967] = 16'hd790;
mem_array[32966] = 16'hbb5b;
mem_array[32969] = 16'hdff9;
mem_array[32968] = 16'hbd28;
mem_array[32971] = 16'h5b7d;
mem_array[32970] = 16'hbe01;
mem_array[32973] = 16'hfcd4;
mem_array[32972] = 16'h3e7c;
mem_array[32975] = 16'hbe08;
mem_array[32974] = 16'hbe07;
mem_array[32977] = 16'h18e0;
mem_array[32976] = 16'h3c10;
mem_array[32979] = 16'h6c23;
mem_array[32978] = 16'hbd3c;
mem_array[32981] = 16'ha238;
mem_array[32980] = 16'hbeb7;
mem_array[32983] = 16'h8ab7;
mem_array[32982] = 16'h3e23;
mem_array[32985] = 16'h966f;
mem_array[32984] = 16'h3dc3;
mem_array[32987] = 16'h9a86;
mem_array[32986] = 16'h3e98;
mem_array[32989] = 16'h6a53;
mem_array[32988] = 16'h3e06;
mem_array[32991] = 16'h25ca;
mem_array[32990] = 16'hbe62;
mem_array[32993] = 16'h5199;
mem_array[32992] = 16'h3e32;
mem_array[32995] = 16'h0b06;
mem_array[32994] = 16'h3e60;
mem_array[32997] = 16'h9a96;
mem_array[32996] = 16'h3e25;
mem_array[32999] = 16'h9772;
mem_array[32998] = 16'hbd40;
mem_array[33001] = 16'h25bc;
mem_array[33000] = 16'hbf81;
mem_array[33003] = 16'h7581;
mem_array[33002] = 16'h3e2c;
mem_array[33005] = 16'h3387;
mem_array[33004] = 16'h3dd0;
mem_array[33007] = 16'h330c;
mem_array[33006] = 16'hbda0;
mem_array[33009] = 16'h0d84;
mem_array[33008] = 16'hbf43;
mem_array[33011] = 16'hbf63;
mem_array[33010] = 16'h3d96;
mem_array[33013] = 16'h4725;
mem_array[33012] = 16'h3e9e;
mem_array[33015] = 16'hca00;
mem_array[33014] = 16'hbe4d;
mem_array[33017] = 16'ha14e;
mem_array[33016] = 16'h3c54;
mem_array[33019] = 16'h4e0f;
mem_array[33018] = 16'h3e64;
mem_array[33021] = 16'h357e;
mem_array[33020] = 16'h3c89;
mem_array[33023] = 16'h9f13;
mem_array[33022] = 16'hbd7f;
mem_array[33025] = 16'h27f1;
mem_array[33024] = 16'hbdeb;
mem_array[33027] = 16'hb76d;
mem_array[33026] = 16'h3e65;
mem_array[33029] = 16'hd837;
mem_array[33028] = 16'h3e18;
mem_array[33031] = 16'hd20a;
mem_array[33030] = 16'hbe95;
mem_array[33033] = 16'h4b8f;
mem_array[33032] = 16'h3f1c;
mem_array[33035] = 16'h5235;
mem_array[33034] = 16'hbdeb;
mem_array[33037] = 16'h3022;
mem_array[33036] = 16'hbee1;
mem_array[33039] = 16'hf100;
mem_array[33038] = 16'h3e4e;
mem_array[33041] = 16'h897d;
mem_array[33040] = 16'hbf0c;
mem_array[33043] = 16'hb2cf;
mem_array[33042] = 16'h3da9;
mem_array[33045] = 16'h12f9;
mem_array[33044] = 16'h3ebc;
mem_array[33047] = 16'h509f;
mem_array[33046] = 16'h3e6f;
mem_array[33049] = 16'hb7f4;
mem_array[33048] = 16'h3e02;
mem_array[33051] = 16'h8124;
mem_array[33050] = 16'hbf2d;
mem_array[33053] = 16'h9cda;
mem_array[33052] = 16'h3e98;
mem_array[33055] = 16'h9385;
mem_array[33054] = 16'h3e92;
mem_array[33057] = 16'hcb82;
mem_array[33056] = 16'h3dea;
mem_array[33059] = 16'hc42a;
mem_array[33058] = 16'hbe4b;
mem_array[33061] = 16'hf55f;
mem_array[33060] = 16'h3e88;
mem_array[33063] = 16'hafd3;
mem_array[33062] = 16'h3d1f;
mem_array[33065] = 16'hd581;
mem_array[33064] = 16'h3e78;
mem_array[33067] = 16'h4245;
mem_array[33066] = 16'hbdf1;
mem_array[33069] = 16'h0314;
mem_array[33068] = 16'hbec4;
mem_array[33071] = 16'hfc73;
mem_array[33070] = 16'hbe3e;
mem_array[33073] = 16'h0fd2;
mem_array[33072] = 16'h3ec3;
mem_array[33075] = 16'hf5a5;
mem_array[33074] = 16'hbec3;
mem_array[33077] = 16'h9abb;
mem_array[33076] = 16'h3dd3;
mem_array[33079] = 16'h41ad;
mem_array[33078] = 16'h3e2b;
mem_array[33081] = 16'hf67e;
mem_array[33080] = 16'h3d27;
mem_array[33083] = 16'h8278;
mem_array[33082] = 16'h3d16;
mem_array[33085] = 16'h6668;
mem_array[33084] = 16'h3df2;
mem_array[33087] = 16'h60b4;
mem_array[33086] = 16'h3d3f;
mem_array[33089] = 16'hc9f6;
mem_array[33088] = 16'h3d21;
mem_array[33091] = 16'h44c7;
mem_array[33090] = 16'hbe1a;
mem_array[33093] = 16'hca6a;
mem_array[33092] = 16'h3df5;
mem_array[33095] = 16'h6a71;
mem_array[33094] = 16'hbbbe;
mem_array[33097] = 16'hfab2;
mem_array[33096] = 16'h3e42;
mem_array[33099] = 16'h29f1;
mem_array[33098] = 16'hbc81;
mem_array[33101] = 16'h0ca7;
mem_array[33100] = 16'hbf59;
mem_array[33103] = 16'hc27c;
mem_array[33102] = 16'h3c54;
mem_array[33105] = 16'h397e;
mem_array[33104] = 16'hbe56;
mem_array[33107] = 16'hb4b4;
mem_array[33106] = 16'h3e3a;
mem_array[33109] = 16'he415;
mem_array[33108] = 16'h3d5b;
mem_array[33111] = 16'h1d1b;
mem_array[33110] = 16'h3e74;
mem_array[33113] = 16'hcd5d;
mem_array[33112] = 16'h3eb1;
mem_array[33115] = 16'he16f;
mem_array[33114] = 16'h3d87;
mem_array[33117] = 16'h8ce6;
mem_array[33116] = 16'hbd1c;
mem_array[33119] = 16'h9334;
mem_array[33118] = 16'h3d65;
mem_array[33121] = 16'h82bd;
mem_array[33120] = 16'hbee6;
mem_array[33123] = 16'h872c;
mem_array[33122] = 16'h3db0;
mem_array[33125] = 16'hfd8a;
mem_array[33124] = 16'h3cc0;
mem_array[33127] = 16'h5e62;
mem_array[33126] = 16'h3d7e;
mem_array[33129] = 16'hd52f;
mem_array[33128] = 16'hbdd4;
mem_array[33131] = 16'h3fe7;
mem_array[33130] = 16'h3e03;
mem_array[33133] = 16'hd383;
mem_array[33132] = 16'h3e38;
mem_array[33135] = 16'h7f34;
mem_array[33134] = 16'hbeca;
mem_array[33137] = 16'h5125;
mem_array[33136] = 16'hbd40;
mem_array[33139] = 16'h16cd;
mem_array[33138] = 16'hbe83;
mem_array[33141] = 16'h389c;
mem_array[33140] = 16'hbde7;
mem_array[33143] = 16'hdf6e;
mem_array[33142] = 16'hbd1d;
mem_array[33145] = 16'h22e1;
mem_array[33144] = 16'h3e94;
mem_array[33147] = 16'h5793;
mem_array[33146] = 16'h3d8e;
mem_array[33149] = 16'h02b3;
mem_array[33148] = 16'hbe3a;
mem_array[33151] = 16'h2c3c;
mem_array[33150] = 16'hbe6c;
mem_array[33153] = 16'h3f1f;
mem_array[33152] = 16'h3e92;
mem_array[33155] = 16'he24f;
mem_array[33154] = 16'hbd75;
mem_array[33157] = 16'h9e56;
mem_array[33156] = 16'hbe8a;
mem_array[33159] = 16'hd46b;
mem_array[33158] = 16'hbe8f;
mem_array[33161] = 16'h201d;
mem_array[33160] = 16'hbf4e;
mem_array[33163] = 16'h06f2;
mem_array[33162] = 16'h3c81;
mem_array[33165] = 16'h3101;
mem_array[33164] = 16'hbe28;
mem_array[33167] = 16'h39d7;
mem_array[33166] = 16'h3e5e;
mem_array[33169] = 16'h20a2;
mem_array[33168] = 16'h3dc4;
mem_array[33171] = 16'h73cb;
mem_array[33170] = 16'hbe6b;
mem_array[33173] = 16'h549e;
mem_array[33172] = 16'h3d69;
mem_array[33175] = 16'h1ea9;
mem_array[33174] = 16'h3dd2;
mem_array[33177] = 16'h4584;
mem_array[33176] = 16'hbb30;
mem_array[33179] = 16'hc9a5;
mem_array[33178] = 16'hbe03;
mem_array[33181] = 16'h5f67;
mem_array[33180] = 16'h3bd1;
mem_array[33183] = 16'h12a1;
mem_array[33182] = 16'hbeee;
mem_array[33185] = 16'h6260;
mem_array[33184] = 16'hbdfe;
mem_array[33187] = 16'h745e;
mem_array[33186] = 16'h3e8d;
mem_array[33189] = 16'h058b;
mem_array[33188] = 16'h3ddd;
mem_array[33191] = 16'h35de;
mem_array[33190] = 16'h3dff;
mem_array[33193] = 16'h48e3;
mem_array[33192] = 16'h3eba;
mem_array[33195] = 16'h3467;
mem_array[33194] = 16'hbf5e;
mem_array[33197] = 16'h1eec;
mem_array[33196] = 16'h3ef5;
mem_array[33199] = 16'h183f;
mem_array[33198] = 16'h3ec5;
mem_array[33201] = 16'h3b7f;
mem_array[33200] = 16'hbb94;
mem_array[33203] = 16'h6025;
mem_array[33202] = 16'hbcec;
mem_array[33205] = 16'hb7a8;
mem_array[33204] = 16'h3d53;
mem_array[33207] = 16'h6186;
mem_array[33206] = 16'h3e1b;
mem_array[33209] = 16'ha245;
mem_array[33208] = 16'h3d1f;
mem_array[33211] = 16'he227;
mem_array[33210] = 16'hbe5a;
mem_array[33213] = 16'hd427;
mem_array[33212] = 16'h3efb;
mem_array[33215] = 16'h2e8f;
mem_array[33214] = 16'hb8a3;
mem_array[33217] = 16'h039c;
mem_array[33216] = 16'hbebb;
mem_array[33219] = 16'hf2ca;
mem_array[33218] = 16'h3cd6;
mem_array[33221] = 16'h5aa6;
mem_array[33220] = 16'hbf89;
mem_array[33223] = 16'hdca8;
mem_array[33222] = 16'h3dd1;
mem_array[33225] = 16'h5f4b;
mem_array[33224] = 16'hbe4e;
mem_array[33227] = 16'hdcf6;
mem_array[33226] = 16'h3e57;
mem_array[33229] = 16'he733;
mem_array[33228] = 16'h3e9e;
mem_array[33231] = 16'hd079;
mem_array[33230] = 16'hbf55;
mem_array[33233] = 16'h1eb7;
mem_array[33232] = 16'h3da1;
mem_array[33235] = 16'h2676;
mem_array[33234] = 16'hbec9;
mem_array[33237] = 16'haf9e;
mem_array[33236] = 16'h3d8b;
mem_array[33239] = 16'h6ea7;
mem_array[33238] = 16'h3e1a;
mem_array[33241] = 16'h374b;
mem_array[33240] = 16'hbee6;
mem_array[33243] = 16'h2834;
mem_array[33242] = 16'hbe88;
mem_array[33245] = 16'hb367;
mem_array[33244] = 16'hbe4a;
mem_array[33247] = 16'h0485;
mem_array[33246] = 16'h3f14;
mem_array[33249] = 16'h2487;
mem_array[33248] = 16'h3e00;
mem_array[33251] = 16'h0976;
mem_array[33250] = 16'h3eb9;
mem_array[33253] = 16'h4d85;
mem_array[33252] = 16'h3eaf;
mem_array[33255] = 16'h16f5;
mem_array[33254] = 16'hbf41;
mem_array[33257] = 16'hce3f;
mem_array[33256] = 16'h3f5d;
mem_array[33259] = 16'h1588;
mem_array[33258] = 16'hbdb9;
mem_array[33261] = 16'hc425;
mem_array[33260] = 16'h3d24;
mem_array[33263] = 16'h81af;
mem_array[33262] = 16'hbba2;
mem_array[33265] = 16'h855d;
mem_array[33264] = 16'h3d4f;
mem_array[33267] = 16'h24f3;
mem_array[33266] = 16'h3c9e;
mem_array[33269] = 16'h17fe;
mem_array[33268] = 16'hbe8b;
mem_array[33271] = 16'h72bb;
mem_array[33270] = 16'hbdba;
mem_array[33273] = 16'hd077;
mem_array[33272] = 16'h3eaa;
mem_array[33275] = 16'h24ed;
mem_array[33274] = 16'h3e9e;
mem_array[33277] = 16'hf4bb;
mem_array[33276] = 16'hbf05;
mem_array[33279] = 16'hc156;
mem_array[33278] = 16'hbf1f;
mem_array[33281] = 16'h77bc;
mem_array[33280] = 16'hc00f;
mem_array[33283] = 16'h1e1c;
mem_array[33282] = 16'hbc13;
mem_array[33285] = 16'h6127;
mem_array[33284] = 16'h3e88;
mem_array[33287] = 16'h1367;
mem_array[33286] = 16'h3e39;
mem_array[33289] = 16'h728c;
mem_array[33288] = 16'h3e6d;
mem_array[33291] = 16'h2d60;
mem_array[33290] = 16'hbf7f;
mem_array[33293] = 16'h92db;
mem_array[33292] = 16'h3e7e;
mem_array[33295] = 16'h970a;
mem_array[33294] = 16'hbe2c;
mem_array[33297] = 16'h3b20;
mem_array[33296] = 16'h3d50;
mem_array[33299] = 16'hc292;
mem_array[33298] = 16'hbf17;
mem_array[33301] = 16'heb24;
mem_array[33300] = 16'hbee5;
mem_array[33303] = 16'hd742;
mem_array[33302] = 16'hbf8b;
mem_array[33305] = 16'h44db;
mem_array[33304] = 16'hbeaa;
mem_array[33307] = 16'h955b;
mem_array[33306] = 16'hbe09;
mem_array[33309] = 16'h73e8;
mem_array[33308] = 16'hbec5;
mem_array[33311] = 16'haadd;
mem_array[33310] = 16'h3eb6;
mem_array[33313] = 16'hebce;
mem_array[33312] = 16'h3ec4;
mem_array[33315] = 16'he8ba;
mem_array[33314] = 16'h3d67;
mem_array[33317] = 16'h8a3a;
mem_array[33316] = 16'h3f02;
mem_array[33319] = 16'hc4ce;
mem_array[33318] = 16'h3e28;
mem_array[33321] = 16'hd904;
mem_array[33320] = 16'hbdff;
mem_array[33323] = 16'h5138;
mem_array[33322] = 16'hbd4e;
mem_array[33325] = 16'h1d17;
mem_array[33324] = 16'hbe81;
mem_array[33327] = 16'h4490;
mem_array[33326] = 16'hbe82;
mem_array[33329] = 16'h56c8;
mem_array[33328] = 16'hbdf3;
mem_array[33331] = 16'hd1c7;
mem_array[33330] = 16'hbdbe;
mem_array[33333] = 16'h665b;
mem_array[33332] = 16'h3d5c;
mem_array[33335] = 16'h1ebf;
mem_array[33334] = 16'h3e45;
mem_array[33337] = 16'h053c;
mem_array[33336] = 16'hbf14;
mem_array[33339] = 16'h7fab;
mem_array[33338] = 16'h3dc1;
mem_array[33341] = 16'hff21;
mem_array[33340] = 16'hbf9f;
mem_array[33343] = 16'h4b86;
mem_array[33342] = 16'h3dae;
mem_array[33345] = 16'ha085;
mem_array[33344] = 16'h3e8e;
mem_array[33347] = 16'hf677;
mem_array[33346] = 16'hbe0e;
mem_array[33349] = 16'h96cb;
mem_array[33348] = 16'h3c26;
mem_array[33351] = 16'h1a2d;
mem_array[33350] = 16'hbd87;
mem_array[33353] = 16'h1f8f;
mem_array[33352] = 16'h3e53;
mem_array[33355] = 16'he4e1;
mem_array[33354] = 16'h3ead;
mem_array[33357] = 16'h0678;
mem_array[33356] = 16'h3e96;
mem_array[33359] = 16'h738d;
mem_array[33358] = 16'hbe7f;
mem_array[33361] = 16'hb801;
mem_array[33360] = 16'hbc9f;
mem_array[33363] = 16'h9ee4;
mem_array[33362] = 16'hbf94;
mem_array[33365] = 16'had69;
mem_array[33364] = 16'hbf05;
mem_array[33367] = 16'h63b5;
mem_array[33366] = 16'hbdf9;
mem_array[33369] = 16'h61e6;
mem_array[33368] = 16'hbf34;
mem_array[33371] = 16'hb2f2;
mem_array[33370] = 16'h3f9d;
mem_array[33373] = 16'h9d78;
mem_array[33372] = 16'h3cbc;
mem_array[33375] = 16'heb78;
mem_array[33374] = 16'h3ed7;
mem_array[33377] = 16'h414a;
mem_array[33376] = 16'h3e02;
mem_array[33379] = 16'h3aa9;
mem_array[33378] = 16'hbede;
mem_array[33381] = 16'hf955;
mem_array[33380] = 16'h3d1b;
mem_array[33383] = 16'hbda4;
mem_array[33382] = 16'hbc77;
mem_array[33385] = 16'h60f0;
mem_array[33384] = 16'hbe89;
mem_array[33387] = 16'hb089;
mem_array[33386] = 16'hbeac;
mem_array[33389] = 16'heb2b;
mem_array[33388] = 16'h3e9d;
mem_array[33391] = 16'hb358;
mem_array[33390] = 16'hbd95;
mem_array[33393] = 16'hf85c;
mem_array[33392] = 16'h3f35;
mem_array[33395] = 16'h919d;
mem_array[33394] = 16'h3ea7;
mem_array[33397] = 16'hb1d1;
mem_array[33396] = 16'hbf4a;
mem_array[33399] = 16'h39b7;
mem_array[33398] = 16'hbe8b;
mem_array[33401] = 16'hb6d3;
mem_array[33400] = 16'hbf57;
mem_array[33403] = 16'h750f;
mem_array[33402] = 16'h3de3;
mem_array[33405] = 16'hc19c;
mem_array[33404] = 16'hbfbf;
mem_array[33407] = 16'h97bd;
mem_array[33406] = 16'hbcb5;
mem_array[33409] = 16'h174c;
mem_array[33408] = 16'hbf1b;
mem_array[33411] = 16'hb946;
mem_array[33410] = 16'h3e23;
mem_array[33413] = 16'hf664;
mem_array[33412] = 16'h3de6;
mem_array[33415] = 16'h012b;
mem_array[33414] = 16'hbf12;
mem_array[33417] = 16'h69cb;
mem_array[33416] = 16'h3eea;
mem_array[33419] = 16'h78f4;
mem_array[33418] = 16'hbdcb;
mem_array[33421] = 16'h9055;
mem_array[33420] = 16'h3f62;
mem_array[33423] = 16'hdc14;
mem_array[33422] = 16'hbe4e;
mem_array[33425] = 16'hff5a;
mem_array[33424] = 16'h3f52;
mem_array[33427] = 16'h9791;
mem_array[33426] = 16'hbf3d;
mem_array[33429] = 16'ha1df;
mem_array[33428] = 16'hbc19;
mem_array[33431] = 16'ha9bb;
mem_array[33430] = 16'h3f64;
mem_array[33433] = 16'h9d8b;
mem_array[33432] = 16'h3c74;
mem_array[33435] = 16'h7b9c;
mem_array[33434] = 16'hba4f;
mem_array[33437] = 16'ha758;
mem_array[33436] = 16'h3de7;
mem_array[33439] = 16'hdda3;
mem_array[33438] = 16'hbec1;
mem_array[33441] = 16'h9b06;
mem_array[33440] = 16'hbc43;
mem_array[33443] = 16'hd279;
mem_array[33442] = 16'h3ce6;
mem_array[33445] = 16'h7e97;
mem_array[33444] = 16'h3b12;
mem_array[33447] = 16'h6a2f;
mem_array[33446] = 16'hbe26;
mem_array[33449] = 16'h9914;
mem_array[33448] = 16'h3f54;
mem_array[33451] = 16'h9203;
mem_array[33450] = 16'hbade;
mem_array[33453] = 16'h3ab2;
mem_array[33452] = 16'h3f05;
mem_array[33455] = 16'heca3;
mem_array[33454] = 16'hbf83;
mem_array[33457] = 16'h12f2;
mem_array[33456] = 16'h3e6e;
mem_array[33459] = 16'ha65e;
mem_array[33458] = 16'hbf3f;
mem_array[33461] = 16'h6bb4;
mem_array[33460] = 16'hbf51;
mem_array[33463] = 16'h4ea8;
mem_array[33462] = 16'hbec4;
mem_array[33465] = 16'hbac3;
mem_array[33464] = 16'hbe2a;
mem_array[33467] = 16'h7361;
mem_array[33466] = 16'h3db3;
mem_array[33469] = 16'hd754;
mem_array[33468] = 16'hbe93;
mem_array[33471] = 16'hf54f;
mem_array[33470] = 16'h3e04;
mem_array[33473] = 16'h9763;
mem_array[33472] = 16'h3de0;
mem_array[33475] = 16'h17e2;
mem_array[33474] = 16'hbf26;
mem_array[33477] = 16'h365d;
mem_array[33476] = 16'h3e34;
mem_array[33479] = 16'hadbe;
mem_array[33478] = 16'hbe60;
mem_array[33481] = 16'hf172;
mem_array[33480] = 16'h3f15;
mem_array[33483] = 16'ha7b1;
mem_array[33482] = 16'h3d0b;
mem_array[33485] = 16'hc168;
mem_array[33484] = 16'h3fc2;
mem_array[33487] = 16'h13bc;
mem_array[33486] = 16'hbf33;
mem_array[33489] = 16'hae77;
mem_array[33488] = 16'h3b57;
mem_array[33491] = 16'h2d1b;
mem_array[33490] = 16'h3c53;
mem_array[33493] = 16'ha9db;
mem_array[33492] = 16'h3f1c;
mem_array[33495] = 16'h49f6;
mem_array[33494] = 16'h3e78;
mem_array[33497] = 16'hc516;
mem_array[33496] = 16'h3f5d;
mem_array[33499] = 16'h7e6d;
mem_array[33498] = 16'h3e72;
mem_array[33501] = 16'h65eb;
mem_array[33500] = 16'hbd1d;
mem_array[33503] = 16'h4e3a;
mem_array[33502] = 16'h3d9b;
mem_array[33505] = 16'h86a5;
mem_array[33504] = 16'hbece;
mem_array[33507] = 16'hd73b;
mem_array[33506] = 16'h3ee0;
mem_array[33509] = 16'ha04a;
mem_array[33508] = 16'h3e8b;
mem_array[33511] = 16'h0476;
mem_array[33510] = 16'h3d9c;
mem_array[33513] = 16'h38db;
mem_array[33512] = 16'h3fc6;
mem_array[33515] = 16'h292d;
mem_array[33514] = 16'h3d08;
mem_array[33517] = 16'h32fe;
mem_array[33516] = 16'h3d0a;
mem_array[33519] = 16'h35d4;
mem_array[33518] = 16'hbe94;
mem_array[33521] = 16'h7605;
mem_array[33520] = 16'h3efa;
mem_array[33523] = 16'hb044;
mem_array[33522] = 16'hbf20;
mem_array[33525] = 16'hb27b;
mem_array[33524] = 16'hbeb0;
mem_array[33527] = 16'h6f9e;
mem_array[33526] = 16'hbf6e;
mem_array[33529] = 16'hb74f;
mem_array[33528] = 16'h3f70;
mem_array[33531] = 16'h7c56;
mem_array[33530] = 16'h3e89;
mem_array[33533] = 16'ha778;
mem_array[33532] = 16'h3f7b;
mem_array[33535] = 16'h04c4;
mem_array[33534] = 16'h3e7e;
mem_array[33537] = 16'hd0e8;
mem_array[33536] = 16'h3f95;
mem_array[33539] = 16'h72be;
mem_array[33538] = 16'hbf20;
mem_array[33541] = 16'hc770;
mem_array[33540] = 16'h3c0f;
mem_array[33543] = 16'hed34;
mem_array[33542] = 16'hbd40;
mem_array[33545] = 16'h67ad;
mem_array[33544] = 16'hbda9;
mem_array[33547] = 16'h2201;
mem_array[33546] = 16'hbe68;
mem_array[33549] = 16'h0ca3;
mem_array[33548] = 16'hbcca;
mem_array[33551] = 16'he1da;
mem_array[33550] = 16'hbe24;
mem_array[33553] = 16'h6507;
mem_array[33552] = 16'h3f3f;
mem_array[33555] = 16'he811;
mem_array[33554] = 16'h3d6d;
mem_array[33557] = 16'hd47e;
mem_array[33556] = 16'h3d80;
mem_array[33559] = 16'h5e06;
mem_array[33558] = 16'h3e01;
mem_array[33561] = 16'hc549;
mem_array[33560] = 16'h3bee;
mem_array[33563] = 16'he129;
mem_array[33562] = 16'hbccb;
mem_array[33565] = 16'h5c6c;
mem_array[33564] = 16'hbe39;
mem_array[33567] = 16'hef62;
mem_array[33566] = 16'h3f41;
mem_array[33569] = 16'h9f81;
mem_array[33568] = 16'h3c01;
mem_array[33571] = 16'h0070;
mem_array[33570] = 16'hbe86;
mem_array[33573] = 16'h95c4;
mem_array[33572] = 16'h3f4b;
mem_array[33575] = 16'h881a;
mem_array[33574] = 16'h3dae;
mem_array[33577] = 16'hf9ab;
mem_array[33576] = 16'h3c74;
mem_array[33579] = 16'h6a00;
mem_array[33578] = 16'h3b82;
mem_array[33581] = 16'ha1e0;
mem_array[33580] = 16'h3e12;
mem_array[33583] = 16'h8d4a;
mem_array[33582] = 16'hbecf;
mem_array[33585] = 16'h301f;
mem_array[33584] = 16'hbe52;
mem_array[33587] = 16'hb8ec;
mem_array[33586] = 16'hbf3b;
mem_array[33589] = 16'h6f45;
mem_array[33588] = 16'h3ee9;
mem_array[33591] = 16'h4e55;
mem_array[33590] = 16'hbdb0;
mem_array[33593] = 16'hcc93;
mem_array[33592] = 16'h3f52;
mem_array[33595] = 16'hea55;
mem_array[33594] = 16'hbd63;
mem_array[33597] = 16'h033e;
mem_array[33596] = 16'h3d33;
mem_array[33599] = 16'h9ced;
mem_array[33598] = 16'hbed9;
mem_array[33601] = 16'he554;
mem_array[33600] = 16'hbd87;
mem_array[33603] = 16'haf8f;
mem_array[33602] = 16'hbd02;
mem_array[33605] = 16'hbfd5;
mem_array[33604] = 16'hbdae;
mem_array[33607] = 16'h4c7c;
mem_array[33606] = 16'hbd34;
mem_array[33609] = 16'h85f3;
mem_array[33608] = 16'hbdab;
mem_array[33611] = 16'h0697;
mem_array[33610] = 16'hbd8b;
mem_array[33613] = 16'hf9bd;
mem_array[33612] = 16'h3d85;
mem_array[33615] = 16'h7591;
mem_array[33614] = 16'hbbc2;
mem_array[33617] = 16'h8068;
mem_array[33616] = 16'h3d5f;
mem_array[33619] = 16'h7871;
mem_array[33618] = 16'h3cc8;
mem_array[33621] = 16'h74eb;
mem_array[33620] = 16'hbc6c;
mem_array[33623] = 16'h8533;
mem_array[33622] = 16'h3d94;
mem_array[33625] = 16'hc137;
mem_array[33624] = 16'hbcf4;
mem_array[33627] = 16'hb3c1;
mem_array[33626] = 16'hbd9e;
mem_array[33629] = 16'h2590;
mem_array[33628] = 16'hbc82;
mem_array[33631] = 16'h3753;
mem_array[33630] = 16'hbd64;
mem_array[33633] = 16'h4a4a;
mem_array[33632] = 16'hbcab;
mem_array[33635] = 16'h634c;
mem_array[33634] = 16'h3d82;
mem_array[33637] = 16'h2039;
mem_array[33636] = 16'h3b14;
mem_array[33639] = 16'h85d8;
mem_array[33638] = 16'hbc8e;
mem_array[33641] = 16'hf6bd;
mem_array[33640] = 16'h3d9b;
mem_array[33643] = 16'hfe0c;
mem_array[33642] = 16'h3d3b;
mem_array[33645] = 16'h448a;
mem_array[33644] = 16'h3d07;
mem_array[33647] = 16'hf4aa;
mem_array[33646] = 16'hbd90;
mem_array[33649] = 16'hd53f;
mem_array[33648] = 16'h3d4b;
mem_array[33651] = 16'h1deb;
mem_array[33650] = 16'h3c80;
mem_array[33653] = 16'he373;
mem_array[33652] = 16'h3d40;
mem_array[33655] = 16'hc2d5;
mem_array[33654] = 16'h3daa;
mem_array[33657] = 16'hceea;
mem_array[33656] = 16'hbc33;
mem_array[33659] = 16'hb14b;
mem_array[33658] = 16'h3bd6;
mem_array[33661] = 16'haf8b;
mem_array[33660] = 16'hbcae;
mem_array[33663] = 16'h85dc;
mem_array[33662] = 16'hbc06;
mem_array[33665] = 16'hc109;
mem_array[33664] = 16'h3e56;
mem_array[33667] = 16'h96cf;
mem_array[33666] = 16'h3d7a;
mem_array[33669] = 16'h6253;
mem_array[33668] = 16'hbd36;
mem_array[33671] = 16'haad9;
mem_array[33670] = 16'hbe9d;
mem_array[33673] = 16'h9cba;
mem_array[33672] = 16'h3e5f;
mem_array[33675] = 16'h2266;
mem_array[33674] = 16'hbdc3;
mem_array[33677] = 16'h1f6e;
mem_array[33676] = 16'hbba0;
mem_array[33679] = 16'h5a5c;
mem_array[33678] = 16'h3da3;
mem_array[33681] = 16'hf4f3;
mem_array[33680] = 16'hbcdc;
mem_array[33683] = 16'h49c6;
mem_array[33682] = 16'hbd16;
mem_array[33685] = 16'h9932;
mem_array[33684] = 16'hbec1;
mem_array[33687] = 16'h07f6;
mem_array[33686] = 16'h3e8b;
mem_array[33689] = 16'h23d2;
mem_array[33688] = 16'h3e91;
mem_array[33691] = 16'he559;
mem_array[33690] = 16'h3dab;
mem_array[33693] = 16'hf196;
mem_array[33692] = 16'hbcb7;
mem_array[33695] = 16'h5a03;
mem_array[33694] = 16'h3d04;
mem_array[33697] = 16'hd33c;
mem_array[33696] = 16'h3e9c;
mem_array[33699] = 16'h27a8;
mem_array[33698] = 16'h3ce4;
mem_array[33701] = 16'h3d3c;
mem_array[33700] = 16'h3e18;
mem_array[33703] = 16'hba4a;
mem_array[33702] = 16'h3ee8;
mem_array[33705] = 16'hdb48;
mem_array[33704] = 16'h3d26;
mem_array[33707] = 16'hcc49;
mem_array[33706] = 16'hbd89;
mem_array[33709] = 16'h9231;
mem_array[33708] = 16'h3dc4;
mem_array[33711] = 16'h1ac1;
mem_array[33710] = 16'h3d34;
mem_array[33713] = 16'h5acf;
mem_array[33712] = 16'hbcde;
mem_array[33715] = 16'h83c3;
mem_array[33714] = 16'h3d57;
mem_array[33717] = 16'h688b;
mem_array[33716] = 16'h3d32;
mem_array[33719] = 16'ha6ee;
mem_array[33718] = 16'hbe16;
mem_array[33721] = 16'h1064;
mem_array[33720] = 16'h3e18;
mem_array[33723] = 16'hb59c;
mem_array[33722] = 16'h3f5a;
mem_array[33725] = 16'hd0ff;
mem_array[33724] = 16'h3e31;
mem_array[33727] = 16'h01ab;
mem_array[33726] = 16'h3f63;
mem_array[33729] = 16'hf29c;
mem_array[33728] = 16'hbecc;
mem_array[33731] = 16'h5cc4;
mem_array[33730] = 16'h3fbf;
mem_array[33733] = 16'hdc7b;
mem_array[33732] = 16'hbe51;
mem_array[33735] = 16'h5d75;
mem_array[33734] = 16'hbda8;
mem_array[33737] = 16'hb782;
mem_array[33736] = 16'hbe15;
mem_array[33739] = 16'ha426;
mem_array[33738] = 16'hbec7;
mem_array[33741] = 16'h0343;
mem_array[33740] = 16'h3d49;
mem_array[33743] = 16'h92a7;
mem_array[33742] = 16'h3ca3;
mem_array[33745] = 16'hf3f7;
mem_array[33744] = 16'hbedd;
mem_array[33747] = 16'h8269;
mem_array[33746] = 16'h3efa;
mem_array[33749] = 16'h1115;
mem_array[33748] = 16'hbdcf;
mem_array[33751] = 16'h54aa;
mem_array[33750] = 16'h3e2b;
mem_array[33753] = 16'hbefa;
mem_array[33752] = 16'hbdbd;
mem_array[33755] = 16'h5872;
mem_array[33754] = 16'h3f12;
mem_array[33757] = 16'hade3;
mem_array[33756] = 16'h3e31;
mem_array[33759] = 16'h048f;
mem_array[33758] = 16'h3e24;
mem_array[33761] = 16'h3809;
mem_array[33760] = 16'hbf13;
mem_array[33763] = 16'h30b7;
mem_array[33762] = 16'h3f02;
mem_array[33765] = 16'h74ca;
mem_array[33764] = 16'h3cdf;
mem_array[33767] = 16'hfb06;
mem_array[33766] = 16'hbe07;
mem_array[33769] = 16'h9ab5;
mem_array[33768] = 16'hbf1f;
mem_array[33771] = 16'haa2b;
mem_array[33770] = 16'h3f69;
mem_array[33773] = 16'had04;
mem_array[33772] = 16'hbd9e;
mem_array[33775] = 16'hcb41;
mem_array[33774] = 16'h3c42;
mem_array[33777] = 16'h08d4;
mem_array[33776] = 16'hbdaf;
mem_array[33779] = 16'h563d;
mem_array[33778] = 16'h3e3c;
mem_array[33781] = 16'h6027;
mem_array[33780] = 16'hbe29;
mem_array[33783] = 16'h76dc;
mem_array[33782] = 16'hbf55;
mem_array[33785] = 16'hce18;
mem_array[33784] = 16'h3da1;
mem_array[33787] = 16'h5c43;
mem_array[33786] = 16'hbd81;
mem_array[33789] = 16'h504a;
mem_array[33788] = 16'hbeb3;
mem_array[33791] = 16'h3c8c;
mem_array[33790] = 16'h3c65;
mem_array[33793] = 16'h7dd5;
mem_array[33792] = 16'h3d68;
mem_array[33795] = 16'h1946;
mem_array[33794] = 16'h3f29;
mem_array[33797] = 16'hb38e;
mem_array[33796] = 16'h3eac;
mem_array[33799] = 16'h4044;
mem_array[33798] = 16'hbec1;
mem_array[33801] = 16'h6bac;
mem_array[33800] = 16'hbcab;
mem_array[33803] = 16'h7bf5;
mem_array[33802] = 16'h3ce9;
mem_array[33805] = 16'h052c;
mem_array[33804] = 16'h3dbe;
mem_array[33807] = 16'h6210;
mem_array[33806] = 16'h3e10;
mem_array[33809] = 16'ha78d;
mem_array[33808] = 16'h3d29;
mem_array[33811] = 16'h7c1c;
mem_array[33810] = 16'h3d0c;
mem_array[33813] = 16'hea36;
mem_array[33812] = 16'h3de8;
mem_array[33815] = 16'hec67;
mem_array[33814] = 16'h3d01;
mem_array[33817] = 16'hd295;
mem_array[33816] = 16'hbe06;
mem_array[33819] = 16'h73cb;
mem_array[33818] = 16'h3f0a;
mem_array[33821] = 16'h31a0;
mem_array[33820] = 16'hbe5f;
mem_array[33823] = 16'h5b9a;
mem_array[33822] = 16'h3e30;
mem_array[33825] = 16'h534b;
mem_array[33824] = 16'hbebf;
mem_array[33827] = 16'h788e;
mem_array[33826] = 16'hbe86;
mem_array[33829] = 16'h5246;
mem_array[33828] = 16'h3f6f;
mem_array[33831] = 16'h7f9b;
mem_array[33830] = 16'h3ccf;
mem_array[33833] = 16'h0c20;
mem_array[33832] = 16'h3efa;
mem_array[33835] = 16'hda34;
mem_array[33834] = 16'hbe07;
mem_array[33837] = 16'hf956;
mem_array[33836] = 16'hbd19;
mem_array[33839] = 16'h59ad;
mem_array[33838] = 16'h3e6d;
mem_array[33841] = 16'h0251;
mem_array[33840] = 16'h3f18;
mem_array[33843] = 16'he9cb;
mem_array[33842] = 16'hbf1c;
mem_array[33845] = 16'h1949;
mem_array[33844] = 16'hbcf0;
mem_array[33847] = 16'h445d;
mem_array[33846] = 16'hbcdd;
mem_array[33849] = 16'h896f;
mem_array[33848] = 16'hbf5b;
mem_array[33851] = 16'hf8ab;
mem_array[33850] = 16'hbdd4;
mem_array[33853] = 16'hee71;
mem_array[33852] = 16'h3d1c;
mem_array[33855] = 16'h9094;
mem_array[33854] = 16'h3d3a;
mem_array[33857] = 16'ha23c;
mem_array[33856] = 16'h3e40;
mem_array[33859] = 16'hd0e1;
mem_array[33858] = 16'hbf23;
mem_array[33861] = 16'h0b4b;
mem_array[33860] = 16'hbd67;
mem_array[33863] = 16'h04e3;
mem_array[33862] = 16'hbd06;
mem_array[33865] = 16'hea48;
mem_array[33864] = 16'h3f00;
mem_array[33867] = 16'h98ce;
mem_array[33866] = 16'h3aff;
mem_array[33869] = 16'h6b1c;
mem_array[33868] = 16'hbd45;
mem_array[33871] = 16'h6f08;
mem_array[33870] = 16'hbe11;
mem_array[33873] = 16'haced;
mem_array[33872] = 16'hbcd4;
mem_array[33875] = 16'hf198;
mem_array[33874] = 16'hbf6a;
mem_array[33877] = 16'hd2aa;
mem_array[33876] = 16'hbfcc;
mem_array[33879] = 16'hc83f;
mem_array[33878] = 16'h3ceb;
mem_array[33881] = 16'h8fa2;
mem_array[33880] = 16'h3ea5;
mem_array[33883] = 16'hc28e;
mem_array[33882] = 16'hbe24;
mem_array[33885] = 16'hc9e9;
mem_array[33884] = 16'hbf6d;
mem_array[33887] = 16'h609c;
mem_array[33886] = 16'hb933;
mem_array[33889] = 16'h749c;
mem_array[33888] = 16'h3e95;
mem_array[33891] = 16'h3991;
mem_array[33890] = 16'hbeaf;
mem_array[33893] = 16'hb35c;
mem_array[33892] = 16'hbb91;
mem_array[33895] = 16'he705;
mem_array[33894] = 16'h3edc;
mem_array[33897] = 16'h4d81;
mem_array[33896] = 16'hbd50;
mem_array[33899] = 16'h5b8a;
mem_array[33898] = 16'hbe4e;
mem_array[33901] = 16'h7ca7;
mem_array[33900] = 16'hbea9;
mem_array[33903] = 16'h62c9;
mem_array[33902] = 16'hbeaa;
mem_array[33905] = 16'h45df;
mem_array[33904] = 16'h3ead;
mem_array[33907] = 16'h8dda;
mem_array[33906] = 16'h3dcc;
mem_array[33909] = 16'h44bb;
mem_array[33908] = 16'hbf00;
mem_array[33911] = 16'he535;
mem_array[33910] = 16'h3e20;
mem_array[33913] = 16'hbaa6;
mem_array[33912] = 16'h3e24;
mem_array[33915] = 16'hf22d;
mem_array[33914] = 16'hbe1e;
mem_array[33917] = 16'h1626;
mem_array[33916] = 16'h3def;
mem_array[33919] = 16'h874f;
mem_array[33918] = 16'hbfae;
mem_array[33921] = 16'h31d3;
mem_array[33920] = 16'h39ec;
mem_array[33923] = 16'h9efd;
mem_array[33922] = 16'hbd3e;
mem_array[33925] = 16'h7a77;
mem_array[33924] = 16'h3e30;
mem_array[33927] = 16'he951;
mem_array[33926] = 16'h3eb1;
mem_array[33929] = 16'h7612;
mem_array[33928] = 16'h3e35;
mem_array[33931] = 16'h7973;
mem_array[33930] = 16'hbe49;
mem_array[33933] = 16'ha404;
mem_array[33932] = 16'h3eab;
mem_array[33935] = 16'hcdd1;
mem_array[33934] = 16'hbea9;
mem_array[33937] = 16'h458a;
mem_array[33936] = 16'hbef5;
mem_array[33939] = 16'h553a;
mem_array[33938] = 16'hbd44;
mem_array[33941] = 16'h5709;
mem_array[33940] = 16'h3df6;
mem_array[33943] = 16'hbc41;
mem_array[33942] = 16'hbe4a;
mem_array[33945] = 16'hde69;
mem_array[33944] = 16'hbf2b;
mem_array[33947] = 16'h4271;
mem_array[33946] = 16'h3d89;
mem_array[33949] = 16'h0706;
mem_array[33948] = 16'h3eef;
mem_array[33951] = 16'h4beb;
mem_array[33950] = 16'hbf0a;
mem_array[33953] = 16'h7361;
mem_array[33952] = 16'h3da1;
mem_array[33955] = 16'hfdc6;
mem_array[33954] = 16'h3e6d;
mem_array[33957] = 16'h2c0e;
mem_array[33956] = 16'h3ef2;
mem_array[33959] = 16'hf4d3;
mem_array[33958] = 16'hbf37;
mem_array[33961] = 16'h4051;
mem_array[33960] = 16'hbc39;
mem_array[33963] = 16'he80b;
mem_array[33962] = 16'hbf2a;
mem_array[33965] = 16'h6011;
mem_array[33964] = 16'h3e3d;
mem_array[33967] = 16'h3f34;
mem_array[33966] = 16'hbb96;
mem_array[33969] = 16'h00c8;
mem_array[33968] = 16'hbf1f;
mem_array[33971] = 16'h1d19;
mem_array[33970] = 16'hbe3e;
mem_array[33973] = 16'h0b11;
mem_array[33972] = 16'h3c58;
mem_array[33975] = 16'h046e;
mem_array[33974] = 16'hbddf;
mem_array[33977] = 16'h8c44;
mem_array[33976] = 16'hbd52;
mem_array[33979] = 16'h7014;
mem_array[33978] = 16'hbf48;
mem_array[33981] = 16'heac6;
mem_array[33980] = 16'hbd11;
mem_array[33983] = 16'h5210;
mem_array[33982] = 16'hbc80;
mem_array[33985] = 16'h02e8;
mem_array[33984] = 16'hbe58;
mem_array[33987] = 16'h5388;
mem_array[33986] = 16'h3cf8;
mem_array[33989] = 16'hd6a5;
mem_array[33988] = 16'h3ddc;
mem_array[33991] = 16'h32f8;
mem_array[33990] = 16'hbc60;
mem_array[33993] = 16'h7f9c;
mem_array[33992] = 16'hbead;
mem_array[33995] = 16'hfdf8;
mem_array[33994] = 16'hbec6;
mem_array[33997] = 16'h5342;
mem_array[33996] = 16'hbeab;
mem_array[33999] = 16'ha89d;
mem_array[33998] = 16'h3e00;
mem_array[34001] = 16'hf3d1;
mem_array[34000] = 16'hbffe;
mem_array[34003] = 16'h32e6;
mem_array[34002] = 16'h3e9f;
mem_array[34005] = 16'hc060;
mem_array[34004] = 16'h3e33;
mem_array[34007] = 16'he705;
mem_array[34006] = 16'hbd67;
mem_array[34009] = 16'hf492;
mem_array[34008] = 16'h3df3;
mem_array[34011] = 16'hd326;
mem_array[34010] = 16'h3f18;
mem_array[34013] = 16'h5b74;
mem_array[34012] = 16'h3e7a;
mem_array[34015] = 16'h4985;
mem_array[34014] = 16'h3ee8;
mem_array[34017] = 16'h6139;
mem_array[34016] = 16'hbed0;
mem_array[34019] = 16'h86ed;
mem_array[34018] = 16'h3c0c;
mem_array[34021] = 16'h772e;
mem_array[34020] = 16'h3e01;
mem_array[34023] = 16'hd5b1;
mem_array[34022] = 16'hbf63;
mem_array[34025] = 16'h66cf;
mem_array[34024] = 16'h3dbb;
mem_array[34027] = 16'hbeac;
mem_array[34026] = 16'h3df0;
mem_array[34029] = 16'h0451;
mem_array[34028] = 16'hbe3d;
mem_array[34031] = 16'hbd46;
mem_array[34030] = 16'hbe17;
mem_array[34033] = 16'h4ca2;
mem_array[34032] = 16'h3dbb;
mem_array[34035] = 16'h324d;
mem_array[34034] = 16'hbde3;
mem_array[34037] = 16'h59f6;
mem_array[34036] = 16'hbddd;
mem_array[34039] = 16'h1eb9;
mem_array[34038] = 16'hbf21;
mem_array[34041] = 16'h791c;
mem_array[34040] = 16'h3c61;
mem_array[34043] = 16'h677a;
mem_array[34042] = 16'hbdca;
mem_array[34045] = 16'h01e6;
mem_array[34044] = 16'h3bcc;
mem_array[34047] = 16'h8090;
mem_array[34046] = 16'h3e89;
mem_array[34049] = 16'hd305;
mem_array[34048] = 16'h3e25;
mem_array[34051] = 16'hd2a8;
mem_array[34050] = 16'h3d0b;
mem_array[34053] = 16'hfc18;
mem_array[34052] = 16'h3e73;
mem_array[34055] = 16'ha944;
mem_array[34054] = 16'hbeab;
mem_array[34057] = 16'hdd5e;
mem_array[34056] = 16'hbf25;
mem_array[34059] = 16'h6562;
mem_array[34058] = 16'h3e3a;
mem_array[34061] = 16'hd198;
mem_array[34060] = 16'hbfbc;
mem_array[34063] = 16'h60e7;
mem_array[34062] = 16'h3dbf;
mem_array[34065] = 16'h3771;
mem_array[34064] = 16'hbc76;
mem_array[34067] = 16'h2f4a;
mem_array[34066] = 16'h3c51;
mem_array[34069] = 16'hd25c;
mem_array[34068] = 16'hbdbb;
mem_array[34071] = 16'h2aee;
mem_array[34070] = 16'h3f40;
mem_array[34073] = 16'h4e75;
mem_array[34072] = 16'h3e9d;
mem_array[34075] = 16'h7f57;
mem_array[34074] = 16'h3e61;
mem_array[34077] = 16'h65ce;
mem_array[34076] = 16'hbe21;
mem_array[34079] = 16'hb66a;
mem_array[34078] = 16'hbd85;
mem_array[34081] = 16'h1e9c;
mem_array[34080] = 16'h3e08;
mem_array[34083] = 16'h5486;
mem_array[34082] = 16'hbf75;
mem_array[34085] = 16'h2088;
mem_array[34084] = 16'h3ea7;
mem_array[34087] = 16'h0e2c;
mem_array[34086] = 16'hbc42;
mem_array[34089] = 16'h66df;
mem_array[34088] = 16'h3e3f;
mem_array[34091] = 16'hf813;
mem_array[34090] = 16'h3ddd;
mem_array[34093] = 16'h1102;
mem_array[34092] = 16'h3c5c;
mem_array[34095] = 16'hf06a;
mem_array[34094] = 16'hb900;
mem_array[34097] = 16'ha59c;
mem_array[34096] = 16'hbe73;
mem_array[34099] = 16'h7b1a;
mem_array[34098] = 16'hbef4;
mem_array[34101] = 16'h71c0;
mem_array[34100] = 16'h3c6f;
mem_array[34103] = 16'h5fc5;
mem_array[34102] = 16'h3d1d;
mem_array[34105] = 16'h45af;
mem_array[34104] = 16'h3c18;
mem_array[34107] = 16'h8a48;
mem_array[34106] = 16'h3ebb;
mem_array[34109] = 16'h4e2b;
mem_array[34108] = 16'h3f05;
mem_array[34111] = 16'h4004;
mem_array[34110] = 16'hbd21;
mem_array[34113] = 16'h751f;
mem_array[34112] = 16'h3d78;
mem_array[34115] = 16'h7895;
mem_array[34114] = 16'hbef9;
mem_array[34117] = 16'he36f;
mem_array[34116] = 16'hbf8e;
mem_array[34119] = 16'hd189;
mem_array[34118] = 16'hbb3a;
mem_array[34121] = 16'hb5ec;
mem_array[34120] = 16'hbe9f;
mem_array[34123] = 16'h4b74;
mem_array[34122] = 16'h3dd4;
mem_array[34125] = 16'h4586;
mem_array[34124] = 16'h3d03;
mem_array[34127] = 16'h7e23;
mem_array[34126] = 16'h3e39;
mem_array[34129] = 16'hc36e;
mem_array[34128] = 16'h3def;
mem_array[34131] = 16'hd7e5;
mem_array[34130] = 16'hbc0a;
mem_array[34133] = 16'h4f5b;
mem_array[34132] = 16'h3e8e;
mem_array[34135] = 16'h3371;
mem_array[34134] = 16'h3e38;
mem_array[34137] = 16'hacdc;
mem_array[34136] = 16'hbe37;
mem_array[34139] = 16'hecf2;
mem_array[34138] = 16'hbe51;
mem_array[34141] = 16'hdc7f;
mem_array[34140] = 16'h3e18;
mem_array[34143] = 16'h92f2;
mem_array[34142] = 16'hbfba;
mem_array[34145] = 16'h1715;
mem_array[34144] = 16'hbdd4;
mem_array[34147] = 16'h87da;
mem_array[34146] = 16'h3f03;
mem_array[34149] = 16'hae5b;
mem_array[34148] = 16'h3c4b;
mem_array[34151] = 16'h22b6;
mem_array[34150] = 16'h3e9d;
mem_array[34153] = 16'h1c38;
mem_array[34152] = 16'h3d9c;
mem_array[34155] = 16'h5430;
mem_array[34154] = 16'hbbe0;
mem_array[34157] = 16'h3de4;
mem_array[34156] = 16'hbe6e;
mem_array[34159] = 16'h5b8c;
mem_array[34158] = 16'h3ee6;
mem_array[34161] = 16'hcfe8;
mem_array[34160] = 16'hbe0c;
mem_array[34163] = 16'hfbb7;
mem_array[34162] = 16'hbdec;
mem_array[34165] = 16'h9fdb;
mem_array[34164] = 16'h3cea;
mem_array[34167] = 16'h1f42;
mem_array[34166] = 16'h3e93;
mem_array[34169] = 16'hf2ff;
mem_array[34168] = 16'h3dfb;
mem_array[34171] = 16'h0bc4;
mem_array[34170] = 16'hbd9a;
mem_array[34173] = 16'hdd36;
mem_array[34172] = 16'h3db8;
mem_array[34175] = 16'h39e9;
mem_array[34174] = 16'hbf50;
mem_array[34177] = 16'h7f28;
mem_array[34176] = 16'hbf44;
mem_array[34179] = 16'h788f;
mem_array[34178] = 16'hbf19;
mem_array[34181] = 16'h4097;
mem_array[34180] = 16'h3f1d;
mem_array[34183] = 16'h325a;
mem_array[34182] = 16'h3cfe;
mem_array[34185] = 16'h51ec;
mem_array[34184] = 16'hbe22;
mem_array[34187] = 16'hda05;
mem_array[34186] = 16'h3e5e;
mem_array[34189] = 16'hf088;
mem_array[34188] = 16'h3dc7;
mem_array[34191] = 16'h3f1a;
mem_array[34190] = 16'hbe88;
mem_array[34193] = 16'h8f37;
mem_array[34192] = 16'h3e42;
mem_array[34195] = 16'ha7dd;
mem_array[34194] = 16'hbd4e;
mem_array[34197] = 16'h1320;
mem_array[34196] = 16'hbe1c;
mem_array[34199] = 16'hd556;
mem_array[34198] = 16'h3d9c;
mem_array[34201] = 16'h5a06;
mem_array[34200] = 16'h3e1d;
mem_array[34203] = 16'h75fb;
mem_array[34202] = 16'hbcb7;
mem_array[34205] = 16'h2bc5;
mem_array[34204] = 16'h3dab;
mem_array[34207] = 16'hc993;
mem_array[34206] = 16'h3ee8;
mem_array[34209] = 16'h6c9d;
mem_array[34208] = 16'h3d68;
mem_array[34211] = 16'h08b2;
mem_array[34210] = 16'h3ec7;
mem_array[34213] = 16'h99a3;
mem_array[34212] = 16'h3d23;
mem_array[34215] = 16'h85ba;
mem_array[34214] = 16'h3d36;
mem_array[34217] = 16'hb18e;
mem_array[34216] = 16'h3e44;
mem_array[34219] = 16'hede0;
mem_array[34218] = 16'hbe65;
mem_array[34221] = 16'h89a3;
mem_array[34220] = 16'hbdd6;
mem_array[34223] = 16'h721a;
mem_array[34222] = 16'hbd02;
mem_array[34225] = 16'hfd6c;
mem_array[34224] = 16'h3ede;
mem_array[34227] = 16'hb3c4;
mem_array[34226] = 16'h3df7;
mem_array[34229] = 16'hc089;
mem_array[34228] = 16'h3dda;
mem_array[34231] = 16'h1f49;
mem_array[34230] = 16'h3c4a;
mem_array[34233] = 16'hf2ae;
mem_array[34232] = 16'h3e23;
mem_array[34235] = 16'h488a;
mem_array[34234] = 16'hbe69;
mem_array[34237] = 16'h2a0d;
mem_array[34236] = 16'hbf81;
mem_array[34239] = 16'h875f;
mem_array[34238] = 16'hbed1;
mem_array[34241] = 16'h160d;
mem_array[34240] = 16'hbb96;
mem_array[34243] = 16'h3e9d;
mem_array[34242] = 16'h3dc1;
mem_array[34245] = 16'h5669;
mem_array[34244] = 16'hbc24;
mem_array[34247] = 16'h80d5;
mem_array[34246] = 16'h3e85;
mem_array[34249] = 16'hc2ab;
mem_array[34248] = 16'hbdee;
mem_array[34251] = 16'h1f39;
mem_array[34250] = 16'hbe7d;
mem_array[34253] = 16'h77f8;
mem_array[34252] = 16'h3e41;
mem_array[34255] = 16'he09e;
mem_array[34254] = 16'h3e09;
mem_array[34257] = 16'hac33;
mem_array[34256] = 16'h3e1f;
mem_array[34259] = 16'hb59d;
mem_array[34258] = 16'h3eb0;
mem_array[34261] = 16'h6372;
mem_array[34260] = 16'h3ed9;
mem_array[34263] = 16'h4831;
mem_array[34262] = 16'h3cb9;
mem_array[34265] = 16'h5a48;
mem_array[34264] = 16'h3ed8;
mem_array[34267] = 16'h334c;
mem_array[34266] = 16'h3ed5;
mem_array[34269] = 16'h84ec;
mem_array[34268] = 16'h3e8e;
mem_array[34271] = 16'hf073;
mem_array[34270] = 16'h3e5d;
mem_array[34273] = 16'h3bdb;
mem_array[34272] = 16'hbd47;
mem_array[34275] = 16'h2c7e;
mem_array[34274] = 16'h3dd0;
mem_array[34277] = 16'h788c;
mem_array[34276] = 16'h3e1d;
mem_array[34279] = 16'h726c;
mem_array[34278] = 16'h3c8b;
mem_array[34281] = 16'hdc58;
mem_array[34280] = 16'hbdce;
mem_array[34283] = 16'h2fe1;
mem_array[34282] = 16'h3d39;
mem_array[34285] = 16'h69e4;
mem_array[34284] = 16'h3eea;
mem_array[34287] = 16'h1ca3;
mem_array[34286] = 16'h3e31;
mem_array[34289] = 16'h0fb8;
mem_array[34288] = 16'h3dd9;
mem_array[34291] = 16'hcd5f;
mem_array[34290] = 16'hbd12;
mem_array[34293] = 16'h810d;
mem_array[34292] = 16'h3da7;
mem_array[34295] = 16'h91f8;
mem_array[34294] = 16'hbe96;
mem_array[34297] = 16'h4af2;
mem_array[34296] = 16'hbee5;
mem_array[34299] = 16'hfc27;
mem_array[34298] = 16'hbeaf;
mem_array[34301] = 16'hdb25;
mem_array[34300] = 16'h3ada;
mem_array[34303] = 16'h883f;
mem_array[34302] = 16'h3e9c;
mem_array[34305] = 16'h24b8;
mem_array[34304] = 16'h3ea4;
mem_array[34307] = 16'hf6a8;
mem_array[34306] = 16'h3e95;
mem_array[34309] = 16'hf8b5;
mem_array[34308] = 16'hbe96;
mem_array[34311] = 16'h886c;
mem_array[34310] = 16'hbd15;
mem_array[34313] = 16'h474c;
mem_array[34312] = 16'h3e7a;
mem_array[34315] = 16'h6d25;
mem_array[34314] = 16'h3e3e;
mem_array[34317] = 16'h1a99;
mem_array[34316] = 16'h3dfd;
mem_array[34319] = 16'h034d;
mem_array[34318] = 16'h3de6;
mem_array[34321] = 16'h3027;
mem_array[34320] = 16'h3e96;
mem_array[34323] = 16'hb533;
mem_array[34322] = 16'hbe71;
mem_array[34325] = 16'had33;
mem_array[34324] = 16'h3ea5;
mem_array[34327] = 16'h9cbc;
mem_array[34326] = 16'h3e4c;
mem_array[34329] = 16'hea35;
mem_array[34328] = 16'h3e12;
mem_array[34331] = 16'h5ca9;
mem_array[34330] = 16'h3cbe;
mem_array[34333] = 16'h1b86;
mem_array[34332] = 16'h3cec;
mem_array[34335] = 16'habf1;
mem_array[34334] = 16'hbce2;
mem_array[34337] = 16'h5d78;
mem_array[34336] = 16'h3dec;
mem_array[34339] = 16'hfc2d;
mem_array[34338] = 16'h3ee3;
mem_array[34341] = 16'h6b56;
mem_array[34340] = 16'hbd58;
mem_array[34343] = 16'h06e5;
mem_array[34342] = 16'h3c50;
mem_array[34345] = 16'hd2dc;
mem_array[34344] = 16'h3eb1;
mem_array[34347] = 16'h5243;
mem_array[34346] = 16'hbddf;
mem_array[34349] = 16'h85e5;
mem_array[34348] = 16'h3e05;
mem_array[34351] = 16'h1928;
mem_array[34350] = 16'h3c20;
mem_array[34353] = 16'h6e13;
mem_array[34352] = 16'h3d62;
mem_array[34355] = 16'h8093;
mem_array[34354] = 16'hbd85;
mem_array[34357] = 16'h1bf8;
mem_array[34356] = 16'hbe6b;
mem_array[34359] = 16'hab21;
mem_array[34358] = 16'hbe3f;
mem_array[34361] = 16'hd461;
mem_array[34360] = 16'h3dd4;
mem_array[34363] = 16'h4bd7;
mem_array[34362] = 16'h3dc9;
mem_array[34365] = 16'h2174;
mem_array[34364] = 16'h3e5f;
mem_array[34367] = 16'h1818;
mem_array[34366] = 16'h3ebf;
mem_array[34369] = 16'h9a94;
mem_array[34368] = 16'hbe26;
mem_array[34371] = 16'h7508;
mem_array[34370] = 16'h3c90;
mem_array[34373] = 16'h4435;
mem_array[34372] = 16'h3d2d;
mem_array[34375] = 16'hf132;
mem_array[34374] = 16'h3de8;
mem_array[34377] = 16'h5656;
mem_array[34376] = 16'hbeb9;
mem_array[34379] = 16'hf087;
mem_array[34378] = 16'h3ebd;
mem_array[34381] = 16'h466e;
mem_array[34380] = 16'hbe90;
mem_array[34383] = 16'h7418;
mem_array[34382] = 16'h3e86;
mem_array[34385] = 16'hfdea;
mem_array[34384] = 16'h3e19;
mem_array[34387] = 16'hd3c2;
mem_array[34386] = 16'h3d7e;
mem_array[34389] = 16'hf55e;
mem_array[34388] = 16'hbd90;
mem_array[34391] = 16'hbfa2;
mem_array[34390] = 16'hbd71;
mem_array[34393] = 16'hc8dc;
mem_array[34392] = 16'h3e34;
mem_array[34395] = 16'h0a77;
mem_array[34394] = 16'h3ea8;
mem_array[34397] = 16'hc2ea;
mem_array[34396] = 16'hbe91;
mem_array[34399] = 16'ha5e2;
mem_array[34398] = 16'h3e28;
mem_array[34401] = 16'h33bd;
mem_array[34400] = 16'hbd90;
mem_array[34403] = 16'hc6be;
mem_array[34402] = 16'hbd71;
mem_array[34405] = 16'h22cf;
mem_array[34404] = 16'h3e49;
mem_array[34407] = 16'he3e3;
mem_array[34406] = 16'hbec5;
mem_array[34409] = 16'hbf5c;
mem_array[34408] = 16'h3d73;
mem_array[34411] = 16'h63d7;
mem_array[34410] = 16'h3dbf;
mem_array[34413] = 16'h5ff6;
mem_array[34412] = 16'h3d23;
mem_array[34415] = 16'hdb75;
mem_array[34414] = 16'h3e3a;
mem_array[34417] = 16'h19c6;
mem_array[34416] = 16'hbe58;
mem_array[34419] = 16'h6e8b;
mem_array[34418] = 16'hbe05;
mem_array[34421] = 16'h4e06;
mem_array[34420] = 16'h3d4f;
mem_array[34423] = 16'h5bc8;
mem_array[34422] = 16'h3e98;
mem_array[34425] = 16'hc444;
mem_array[34424] = 16'h3f14;
mem_array[34427] = 16'h8903;
mem_array[34426] = 16'h3e2c;
mem_array[34429] = 16'h6c67;
mem_array[34428] = 16'hbe50;
mem_array[34431] = 16'hd717;
mem_array[34430] = 16'hbea2;
mem_array[34433] = 16'h3142;
mem_array[34432] = 16'hbd0c;
mem_array[34435] = 16'h7043;
mem_array[34434] = 16'h3bc6;
mem_array[34437] = 16'hce58;
mem_array[34436] = 16'hbed8;
mem_array[34439] = 16'h5c43;
mem_array[34438] = 16'h3ee5;
mem_array[34441] = 16'h2544;
mem_array[34440] = 16'hbedf;
mem_array[34443] = 16'h7ad3;
mem_array[34442] = 16'h3eca;
mem_array[34445] = 16'hfc38;
mem_array[34444] = 16'h3cef;
mem_array[34447] = 16'hf161;
mem_array[34446] = 16'hbe30;
mem_array[34449] = 16'h8559;
mem_array[34448] = 16'hbf03;
mem_array[34451] = 16'hcd6e;
mem_array[34450] = 16'h3de6;
mem_array[34453] = 16'h7160;
mem_array[34452] = 16'h3d4b;
mem_array[34455] = 16'h270e;
mem_array[34454] = 16'h3d9a;
mem_array[34457] = 16'h15a3;
mem_array[34456] = 16'hbe83;
mem_array[34459] = 16'h5eae;
mem_array[34458] = 16'h3e32;
mem_array[34461] = 16'hd8fe;
mem_array[34460] = 16'hbcce;
mem_array[34463] = 16'hb1a2;
mem_array[34462] = 16'h3d7c;
mem_array[34465] = 16'hc2a5;
mem_array[34464] = 16'h3e9f;
mem_array[34467] = 16'h6f0f;
mem_array[34466] = 16'hbe0d;
mem_array[34469] = 16'h3df6;
mem_array[34468] = 16'h3e54;
mem_array[34471] = 16'h499a;
mem_array[34470] = 16'hbe41;
mem_array[34473] = 16'h131b;
mem_array[34472] = 16'hbda9;
mem_array[34475] = 16'hc510;
mem_array[34474] = 16'hbdbf;
mem_array[34477] = 16'h9e4f;
mem_array[34476] = 16'hbd49;
mem_array[34479] = 16'h7044;
mem_array[34478] = 16'h3b8c;
mem_array[34481] = 16'hd78c;
mem_array[34480] = 16'h3e6d;
mem_array[34483] = 16'hfbe0;
mem_array[34482] = 16'h3d4c;
mem_array[34485] = 16'h8901;
mem_array[34484] = 16'h3ea0;
mem_array[34487] = 16'h77a3;
mem_array[34486] = 16'hbe1b;
mem_array[34489] = 16'h1721;
mem_array[34488] = 16'hbd7f;
mem_array[34491] = 16'he747;
mem_array[34490] = 16'h3e88;
mem_array[34493] = 16'hdf4a;
mem_array[34492] = 16'h3ccf;
mem_array[34495] = 16'h9e6d;
mem_array[34494] = 16'hbe0e;
mem_array[34497] = 16'h6dc9;
mem_array[34496] = 16'hbf5f;
mem_array[34499] = 16'hb7d5;
mem_array[34498] = 16'h3edc;
mem_array[34501] = 16'hc7bc;
mem_array[34500] = 16'hbf14;
mem_array[34503] = 16'he84d;
mem_array[34502] = 16'hbda8;
mem_array[34505] = 16'h7a8e;
mem_array[34504] = 16'hbca8;
mem_array[34507] = 16'h96ff;
mem_array[34506] = 16'hbdf4;
mem_array[34509] = 16'h97ba;
mem_array[34508] = 16'hbf20;
mem_array[34511] = 16'h61c6;
mem_array[34510] = 16'hbd51;
mem_array[34513] = 16'h8d32;
mem_array[34512] = 16'hbdb8;
mem_array[34515] = 16'h206b;
mem_array[34514] = 16'h3dc9;
mem_array[34517] = 16'h6ec1;
mem_array[34516] = 16'hbed5;
mem_array[34519] = 16'h0b04;
mem_array[34518] = 16'h3cef;
mem_array[34521] = 16'hfe5f;
mem_array[34520] = 16'hbcff;
mem_array[34523] = 16'h9b75;
mem_array[34522] = 16'hbd5c;
mem_array[34525] = 16'hcb03;
mem_array[34524] = 16'hbd2f;
mem_array[34527] = 16'h6bde;
mem_array[34526] = 16'hbd05;
mem_array[34529] = 16'h55e0;
mem_array[34528] = 16'h3e2f;
mem_array[34531] = 16'h02c6;
mem_array[34530] = 16'hbdab;
mem_array[34533] = 16'h797e;
mem_array[34532] = 16'h3e93;
mem_array[34535] = 16'h4156;
mem_array[34534] = 16'h3c64;
mem_array[34537] = 16'h7c4e;
mem_array[34536] = 16'hbec9;
mem_array[34539] = 16'h49d5;
mem_array[34538] = 16'h3e61;
mem_array[34541] = 16'hf3bf;
mem_array[34540] = 16'hbe7d;
mem_array[34543] = 16'h41d0;
mem_array[34542] = 16'h3e5a;
mem_array[34545] = 16'h0c43;
mem_array[34544] = 16'h3ec9;
mem_array[34547] = 16'h67ab;
mem_array[34546] = 16'h3c99;
mem_array[34549] = 16'haad4;
mem_array[34548] = 16'hbdae;
mem_array[34551] = 16'h4178;
mem_array[34550] = 16'h3d48;
mem_array[34553] = 16'hcbdc;
mem_array[34552] = 16'h3eb4;
mem_array[34555] = 16'h507c;
mem_array[34554] = 16'hbd53;
mem_array[34557] = 16'h055b;
mem_array[34556] = 16'hbf3f;
mem_array[34559] = 16'h8d73;
mem_array[34558] = 16'h3e70;
mem_array[34561] = 16'h4ed7;
mem_array[34560] = 16'hbf1a;
mem_array[34563] = 16'h249b;
mem_array[34562] = 16'h3cc2;
mem_array[34565] = 16'h572a;
mem_array[34564] = 16'h3d03;
mem_array[34567] = 16'h1572;
mem_array[34566] = 16'hbdad;
mem_array[34569] = 16'h9be7;
mem_array[34568] = 16'hbf19;
mem_array[34571] = 16'h90d8;
mem_array[34570] = 16'h3d9c;
mem_array[34573] = 16'h3b38;
mem_array[34572] = 16'hbe10;
mem_array[34575] = 16'h191d;
mem_array[34574] = 16'h3c10;
mem_array[34577] = 16'h2f3f;
mem_array[34576] = 16'hbeb1;
mem_array[34579] = 16'h48bc;
mem_array[34578] = 16'h3ea3;
mem_array[34581] = 16'h172f;
mem_array[34580] = 16'hbc5c;
mem_array[34583] = 16'h2372;
mem_array[34582] = 16'hbb6c;
mem_array[34585] = 16'h6149;
mem_array[34584] = 16'hbdd0;
mem_array[34587] = 16'heee8;
mem_array[34586] = 16'h3e71;
mem_array[34589] = 16'hebbb;
mem_array[34588] = 16'h3e83;
mem_array[34591] = 16'hf4ef;
mem_array[34590] = 16'h3daa;
mem_array[34593] = 16'hb5a7;
mem_array[34592] = 16'h3e58;
mem_array[34595] = 16'h52bb;
mem_array[34594] = 16'hbacb;
mem_array[34597] = 16'he9d1;
mem_array[34596] = 16'h3d23;
mem_array[34599] = 16'h50f6;
mem_array[34598] = 16'hbd15;
mem_array[34601] = 16'h9021;
mem_array[34600] = 16'hbd46;
mem_array[34603] = 16'h268f;
mem_array[34602] = 16'h3e2c;
mem_array[34605] = 16'hb9fe;
mem_array[34604] = 16'h3c93;
mem_array[34607] = 16'h45a2;
mem_array[34606] = 16'hbd09;
mem_array[34609] = 16'h3eb8;
mem_array[34608] = 16'hbdb6;
mem_array[34611] = 16'had76;
mem_array[34610] = 16'hbe9b;
mem_array[34613] = 16'h4ceb;
mem_array[34612] = 16'h3e44;
mem_array[34615] = 16'hb1a0;
mem_array[34614] = 16'h3e60;
mem_array[34617] = 16'h2162;
mem_array[34616] = 16'hbedc;
mem_array[34619] = 16'he59f;
mem_array[34618] = 16'h3d88;
mem_array[34621] = 16'h3533;
mem_array[34620] = 16'hbda9;
mem_array[34623] = 16'h9ce3;
mem_array[34622] = 16'hbd90;
mem_array[34625] = 16'h6d9c;
mem_array[34624] = 16'hbced;
mem_array[34627] = 16'h4be8;
mem_array[34626] = 16'h3e44;
mem_array[34629] = 16'ha92e;
mem_array[34628] = 16'hbf72;
mem_array[34631] = 16'h84fe;
mem_array[34630] = 16'h3e9a;
mem_array[34633] = 16'h2569;
mem_array[34632] = 16'hbe65;
mem_array[34635] = 16'hd1c1;
mem_array[34634] = 16'hbe9d;
mem_array[34637] = 16'h4875;
mem_array[34636] = 16'hbf0b;
mem_array[34639] = 16'h45bc;
mem_array[34638] = 16'h3e0b;
mem_array[34641] = 16'h2b38;
mem_array[34640] = 16'hbd58;
mem_array[34643] = 16'h6cf6;
mem_array[34642] = 16'hbde1;
mem_array[34645] = 16'h4e3b;
mem_array[34644] = 16'hbc04;
mem_array[34647] = 16'h80f9;
mem_array[34646] = 16'hbd8b;
mem_array[34649] = 16'h4d75;
mem_array[34648] = 16'hbe02;
mem_array[34651] = 16'h4b7e;
mem_array[34650] = 16'h3d83;
mem_array[34653] = 16'h1833;
mem_array[34652] = 16'h3e8c;
mem_array[34655] = 16'h4abd;
mem_array[34654] = 16'h3c35;
mem_array[34657] = 16'h227a;
mem_array[34656] = 16'hbeed;
mem_array[34659] = 16'h9c72;
mem_array[34658] = 16'h3de2;
mem_array[34661] = 16'hdb94;
mem_array[34660] = 16'hbeb8;
mem_array[34663] = 16'h97f1;
mem_array[34662] = 16'h3dcd;
mem_array[34665] = 16'h3948;
mem_array[34664] = 16'h3d80;
mem_array[34667] = 16'h7354;
mem_array[34666] = 16'hbe32;
mem_array[34669] = 16'h3d8e;
mem_array[34668] = 16'hbe6b;
mem_array[34671] = 16'h92c9;
mem_array[34670] = 16'hbe91;
mem_array[34673] = 16'hdba9;
mem_array[34672] = 16'h3e42;
mem_array[34675] = 16'hfe74;
mem_array[34674] = 16'hbe60;
mem_array[34677] = 16'h3ec7;
mem_array[34676] = 16'hbe23;
mem_array[34679] = 16'hcafc;
mem_array[34678] = 16'hbd74;
mem_array[34681] = 16'h34c2;
mem_array[34680] = 16'hbf2f;
mem_array[34683] = 16'h4084;
mem_array[34682] = 16'hbd34;
mem_array[34685] = 16'hf1be;
mem_array[34684] = 16'hbd4d;
mem_array[34687] = 16'h5949;
mem_array[34686] = 16'hbd7e;
mem_array[34689] = 16'ha93b;
mem_array[34688] = 16'hbf19;
mem_array[34691] = 16'hedf0;
mem_array[34690] = 16'h3e46;
mem_array[34693] = 16'h7f15;
mem_array[34692] = 16'h3d8c;
mem_array[34695] = 16'hf86c;
mem_array[34694] = 16'hbe72;
mem_array[34697] = 16'hc2c6;
mem_array[34696] = 16'hbeb8;
mem_array[34699] = 16'hc5ac;
mem_array[34698] = 16'h3ead;
mem_array[34701] = 16'hdfdf;
mem_array[34700] = 16'hbd04;
mem_array[34703] = 16'h472e;
mem_array[34702] = 16'hbd78;
mem_array[34705] = 16'h5b9e;
mem_array[34704] = 16'h3d0c;
mem_array[34707] = 16'h9e57;
mem_array[34706] = 16'h3dd3;
mem_array[34709] = 16'h7b42;
mem_array[34708] = 16'hbe6b;
mem_array[34711] = 16'hf042;
mem_array[34710] = 16'hbc5e;
mem_array[34713] = 16'hdf4d;
mem_array[34712] = 16'h3d23;
mem_array[34715] = 16'hd6e8;
mem_array[34714] = 16'h3d76;
mem_array[34717] = 16'hb7f9;
mem_array[34716] = 16'hbed5;
mem_array[34719] = 16'h7a75;
mem_array[34718] = 16'h3ee9;
mem_array[34721] = 16'h9b39;
mem_array[34720] = 16'hbe5d;
mem_array[34723] = 16'ha450;
mem_array[34722] = 16'hbc3c;
mem_array[34725] = 16'h68e3;
mem_array[34724] = 16'h3e52;
mem_array[34727] = 16'h7e84;
mem_array[34726] = 16'hbe6f;
mem_array[34729] = 16'h0a78;
mem_array[34728] = 16'h3e83;
mem_array[34731] = 16'h6e49;
mem_array[34730] = 16'hbf9b;
mem_array[34733] = 16'hb350;
mem_array[34732] = 16'h3dce;
mem_array[34735] = 16'h4bd8;
mem_array[34734] = 16'hbd41;
mem_array[34737] = 16'h6b64;
mem_array[34736] = 16'hbe98;
mem_array[34739] = 16'h132d;
mem_array[34738] = 16'h3d94;
mem_array[34741] = 16'h2d39;
mem_array[34740] = 16'hbeb2;
mem_array[34743] = 16'hcc87;
mem_array[34742] = 16'hbe65;
mem_array[34745] = 16'h0649;
mem_array[34744] = 16'h3cc9;
mem_array[34747] = 16'h6f49;
mem_array[34746] = 16'hbe77;
mem_array[34749] = 16'h495d;
mem_array[34748] = 16'hbcb8;
mem_array[34751] = 16'hca8d;
mem_array[34750] = 16'hbe27;
mem_array[34753] = 16'h668b;
mem_array[34752] = 16'hbe04;
mem_array[34755] = 16'hdeb9;
mem_array[34754] = 16'hbecb;
mem_array[34757] = 16'hd78e;
mem_array[34756] = 16'hbeb2;
mem_array[34759] = 16'h7992;
mem_array[34758] = 16'h3db0;
mem_array[34761] = 16'h48d9;
mem_array[34760] = 16'h3ca6;
mem_array[34763] = 16'h29bc;
mem_array[34762] = 16'hbd2c;
mem_array[34765] = 16'haec1;
mem_array[34764] = 16'hbdb1;
mem_array[34767] = 16'hecd5;
mem_array[34766] = 16'h3dfb;
mem_array[34769] = 16'hf55a;
mem_array[34768] = 16'hbcce;
mem_array[34771] = 16'h8498;
mem_array[34770] = 16'hbdbf;
mem_array[34773] = 16'hc961;
mem_array[34772] = 16'hbc39;
mem_array[34775] = 16'h52f6;
mem_array[34774] = 16'h3e36;
mem_array[34777] = 16'h7755;
mem_array[34776] = 16'hbec5;
mem_array[34779] = 16'h9388;
mem_array[34778] = 16'h3e68;
mem_array[34781] = 16'h3748;
mem_array[34780] = 16'hbf0c;
mem_array[34783] = 16'h9e22;
mem_array[34782] = 16'hbe2e;
mem_array[34785] = 16'h13c4;
mem_array[34784] = 16'h3e5c;
mem_array[34787] = 16'h158e;
mem_array[34786] = 16'hbe2b;
mem_array[34789] = 16'ha462;
mem_array[34788] = 16'hbe0f;
mem_array[34791] = 16'hc7c2;
mem_array[34790] = 16'hbf35;
mem_array[34793] = 16'h7d8a;
mem_array[34792] = 16'h3e5c;
mem_array[34795] = 16'h727b;
mem_array[34794] = 16'h3e1f;
mem_array[34797] = 16'hab7b;
mem_array[34796] = 16'hbe59;
mem_array[34799] = 16'h88b4;
mem_array[34798] = 16'h3e22;
mem_array[34801] = 16'he1e1;
mem_array[34800] = 16'hbffc;
mem_array[34803] = 16'hefb7;
mem_array[34802] = 16'hbf07;
mem_array[34805] = 16'hddbb;
mem_array[34804] = 16'h3e34;
mem_array[34807] = 16'h7a52;
mem_array[34806] = 16'hbed3;
mem_array[34809] = 16'h8a9f;
mem_array[34808] = 16'h3de9;
mem_array[34811] = 16'h9348;
mem_array[34810] = 16'hbe53;
mem_array[34813] = 16'h4661;
mem_array[34812] = 16'hbd22;
mem_array[34815] = 16'h21ef;
mem_array[34814] = 16'hbeec;
mem_array[34817] = 16'h6a3a;
mem_array[34816] = 16'h3e3b;
mem_array[34819] = 16'h5d93;
mem_array[34818] = 16'hbe09;
mem_array[34821] = 16'hacf3;
mem_array[34820] = 16'h3c42;
mem_array[34823] = 16'hd7b7;
mem_array[34822] = 16'hbdb8;
mem_array[34825] = 16'h6da1;
mem_array[34824] = 16'hbdb7;
mem_array[34827] = 16'h11fa;
mem_array[34826] = 16'h3d1b;
mem_array[34829] = 16'hc696;
mem_array[34828] = 16'h3eb6;
mem_array[34831] = 16'h6ccc;
mem_array[34830] = 16'h3b65;
mem_array[34833] = 16'h61ed;
mem_array[34832] = 16'hbdfb;
mem_array[34835] = 16'h336d;
mem_array[34834] = 16'h3e26;
mem_array[34837] = 16'h9ea0;
mem_array[34836] = 16'hbf46;
mem_array[34839] = 16'h3d5d;
mem_array[34838] = 16'h3ceb;
mem_array[34841] = 16'h5f70;
mem_array[34840] = 16'hbf93;
mem_array[34843] = 16'hbb67;
mem_array[34842] = 16'h3e20;
mem_array[34845] = 16'hd83a;
mem_array[34844] = 16'hbc9f;
mem_array[34847] = 16'h9c84;
mem_array[34846] = 16'h3a94;
mem_array[34849] = 16'h4b5d;
mem_array[34848] = 16'h3d62;
mem_array[34851] = 16'hb866;
mem_array[34850] = 16'hbfbf;
mem_array[34853] = 16'hb7c5;
mem_array[34852] = 16'h3eed;
mem_array[34855] = 16'h762f;
mem_array[34854] = 16'h3ce9;
mem_array[34857] = 16'h30f6;
mem_array[34856] = 16'hbe34;
mem_array[34859] = 16'he581;
mem_array[34858] = 16'h3da7;
mem_array[34861] = 16'h5fc8;
mem_array[34860] = 16'hbf3a;
mem_array[34863] = 16'h6b6c;
mem_array[34862] = 16'hbf53;
mem_array[34865] = 16'hb4ec;
mem_array[34864] = 16'hbd43;
mem_array[34867] = 16'headc;
mem_array[34866] = 16'h3bb9;
mem_array[34869] = 16'h3711;
mem_array[34868] = 16'h3e19;
mem_array[34871] = 16'hb1d0;
mem_array[34870] = 16'h3ea9;
mem_array[34873] = 16'h2c98;
mem_array[34872] = 16'h3e72;
mem_array[34875] = 16'h306c;
mem_array[34874] = 16'hbf4f;
mem_array[34877] = 16'h98e1;
mem_array[34876] = 16'h3e2f;
mem_array[34879] = 16'h4e1b;
mem_array[34878] = 16'hbca8;
mem_array[34881] = 16'h4906;
mem_array[34880] = 16'h3d3a;
mem_array[34883] = 16'hd230;
mem_array[34882] = 16'hbd10;
mem_array[34885] = 16'h8a1d;
mem_array[34884] = 16'hbdcd;
mem_array[34887] = 16'h3493;
mem_array[34886] = 16'hbeda;
mem_array[34889] = 16'hc6fe;
mem_array[34888] = 16'h3deb;
mem_array[34891] = 16'h1dfa;
mem_array[34890] = 16'h3e06;
mem_array[34893] = 16'h94b1;
mem_array[34892] = 16'hbd7d;
mem_array[34895] = 16'h004c;
mem_array[34894] = 16'hbe0b;
mem_array[34897] = 16'h712a;
mem_array[34896] = 16'hbf23;
mem_array[34899] = 16'hd41c;
mem_array[34898] = 16'h3e30;
mem_array[34901] = 16'had43;
mem_array[34900] = 16'hbf6f;
mem_array[34903] = 16'hf12f;
mem_array[34902] = 16'h3e6f;
mem_array[34905] = 16'heff5;
mem_array[34904] = 16'hbe51;
mem_array[34907] = 16'h3332;
mem_array[34906] = 16'h3e5c;
mem_array[34909] = 16'h679b;
mem_array[34908] = 16'hbd56;
mem_array[34911] = 16'h4824;
mem_array[34910] = 16'hbf97;
mem_array[34913] = 16'h5aec;
mem_array[34912] = 16'h3ed5;
mem_array[34915] = 16'h41d4;
mem_array[34914] = 16'h3cc0;
mem_array[34917] = 16'he085;
mem_array[34916] = 16'hbe93;
mem_array[34919] = 16'hcbb6;
mem_array[34918] = 16'hbe0d;
mem_array[34921] = 16'h829a;
mem_array[34920] = 16'hbf05;
mem_array[34923] = 16'hbe1e;
mem_array[34922] = 16'hbe14;
mem_array[34925] = 16'h660b;
mem_array[34924] = 16'h3e09;
mem_array[34927] = 16'hc29b;
mem_array[34926] = 16'hbdd9;
mem_array[34929] = 16'h1c5e;
mem_array[34928] = 16'h3e4d;
mem_array[34931] = 16'h51bc;
mem_array[34930] = 16'hbd7d;
mem_array[34933] = 16'h0e3b;
mem_array[34932] = 16'h3ecf;
mem_array[34935] = 16'h4815;
mem_array[34934] = 16'hbf05;
mem_array[34937] = 16'h8c13;
mem_array[34936] = 16'h3e8e;
mem_array[34939] = 16'h2071;
mem_array[34938] = 16'hbe99;
mem_array[34941] = 16'h0f8d;
mem_array[34940] = 16'hbc29;
mem_array[34943] = 16'he6bf;
mem_array[34942] = 16'hbd07;
mem_array[34945] = 16'h7c56;
mem_array[34944] = 16'hbe8a;
mem_array[34947] = 16'h7e20;
mem_array[34946] = 16'hbeb3;
mem_array[34949] = 16'h8568;
mem_array[34948] = 16'hbda8;
mem_array[34951] = 16'h0b0e;
mem_array[34950] = 16'h3e4e;
mem_array[34953] = 16'h3658;
mem_array[34952] = 16'h3eaf;
mem_array[34955] = 16'h19b7;
mem_array[34954] = 16'h3d8b;
mem_array[34957] = 16'h58f4;
mem_array[34956] = 16'hbebc;
mem_array[34959] = 16'h7059;
mem_array[34958] = 16'h3dee;
mem_array[34961] = 16'hfc90;
mem_array[34960] = 16'hbf93;
mem_array[34963] = 16'h6588;
mem_array[34962] = 16'hbc8b;
mem_array[34965] = 16'h5ebd;
mem_array[34964] = 16'h3d8b;
mem_array[34967] = 16'hdcd2;
mem_array[34966] = 16'h3e7e;
mem_array[34969] = 16'h1b6a;
mem_array[34968] = 16'hbf18;
mem_array[34971] = 16'h9f5b;
mem_array[34970] = 16'hbecf;
mem_array[34973] = 16'h2209;
mem_array[34972] = 16'h3e9c;
mem_array[34975] = 16'hed52;
mem_array[34974] = 16'h3d8d;
mem_array[34977] = 16'hf2da;
mem_array[34976] = 16'h3dcc;
mem_array[34979] = 16'h5f02;
mem_array[34978] = 16'hbf36;
mem_array[34981] = 16'hc2e2;
mem_array[34980] = 16'h3e71;
mem_array[34983] = 16'h73ac;
mem_array[34982] = 16'hbee5;
mem_array[34985] = 16'h8974;
mem_array[34984] = 16'hbc96;
mem_array[34987] = 16'h2daa;
mem_array[34986] = 16'hbde1;
mem_array[34989] = 16'h5547;
mem_array[34988] = 16'h3ddf;
mem_array[34991] = 16'h76d7;
mem_array[34990] = 16'h3d93;
mem_array[34993] = 16'h3b93;
mem_array[34992] = 16'hbeb0;
mem_array[34995] = 16'h13b3;
mem_array[34994] = 16'hbdcb;
mem_array[34997] = 16'h4311;
mem_array[34996] = 16'h3ecc;
mem_array[34999] = 16'hdf7e;
mem_array[34998] = 16'h3e20;
mem_array[35001] = 16'h33ac;
mem_array[35000] = 16'hbdd7;
mem_array[35003] = 16'h0546;
mem_array[35002] = 16'hbb26;
mem_array[35005] = 16'h8594;
mem_array[35004] = 16'hbefc;
mem_array[35007] = 16'h7c75;
mem_array[35006] = 16'h3d1b;
mem_array[35009] = 16'he663;
mem_array[35008] = 16'h3ed0;
mem_array[35011] = 16'h34d0;
mem_array[35010] = 16'h3e3b;
mem_array[35013] = 16'h2202;
mem_array[35012] = 16'h3e38;
mem_array[35015] = 16'h9e5f;
mem_array[35014] = 16'h3dea;
mem_array[35017] = 16'h07dc;
mem_array[35016] = 16'hbf7e;
mem_array[35019] = 16'ha926;
mem_array[35018] = 16'h3f2f;
mem_array[35021] = 16'h9c9c;
mem_array[35020] = 16'hbe1b;
mem_array[35023] = 16'h847a;
mem_array[35022] = 16'h3e85;
mem_array[35025] = 16'h4490;
mem_array[35024] = 16'h3f80;
mem_array[35027] = 16'h6012;
mem_array[35026] = 16'hbe7f;
mem_array[35029] = 16'h27a7;
mem_array[35028] = 16'hbf14;
mem_array[35031] = 16'hd238;
mem_array[35030] = 16'hbf0c;
mem_array[35033] = 16'h6e78;
mem_array[35032] = 16'h3e87;
mem_array[35035] = 16'h74b0;
mem_array[35034] = 16'h3f41;
mem_array[35037] = 16'h2b65;
mem_array[35036] = 16'hbe66;
mem_array[35039] = 16'h83f8;
mem_array[35038] = 16'hbf49;
mem_array[35041] = 16'h35f2;
mem_array[35040] = 16'h3f16;
mem_array[35043] = 16'h0aa3;
mem_array[35042] = 16'hbeab;
mem_array[35045] = 16'hb638;
mem_array[35044] = 16'hbeba;
mem_array[35047] = 16'hd8d5;
mem_array[35046] = 16'hbd5c;
mem_array[35049] = 16'hbd54;
mem_array[35048] = 16'hbea5;
mem_array[35051] = 16'h11d5;
mem_array[35050] = 16'h3fc2;
mem_array[35053] = 16'hf6d1;
mem_array[35052] = 16'h3d35;
mem_array[35055] = 16'hdc62;
mem_array[35054] = 16'hbbac;
mem_array[35057] = 16'h11fb;
mem_array[35056] = 16'h3e8a;
mem_array[35059] = 16'h72ff;
mem_array[35058] = 16'h3de2;
mem_array[35061] = 16'h1539;
mem_array[35060] = 16'h3cec;
mem_array[35063] = 16'h0889;
mem_array[35062] = 16'h3b4e;
mem_array[35065] = 16'h43fa;
mem_array[35064] = 16'hbe98;
mem_array[35067] = 16'h6081;
mem_array[35066] = 16'h3f16;
mem_array[35069] = 16'hc4df;
mem_array[35068] = 16'h3f2b;
mem_array[35071] = 16'h19a0;
mem_array[35070] = 16'hbf0c;
mem_array[35073] = 16'h00d1;
mem_array[35072] = 16'h3edc;
mem_array[35075] = 16'h5b46;
mem_array[35074] = 16'hbe3e;
mem_array[35077] = 16'h39a4;
mem_array[35076] = 16'hbda2;
mem_array[35079] = 16'h3a73;
mem_array[35078] = 16'h3f01;
mem_array[35081] = 16'hba1b;
mem_array[35080] = 16'hbee1;
mem_array[35083] = 16'h83c1;
mem_array[35082] = 16'hbe3c;
mem_array[35085] = 16'h5502;
mem_array[35084] = 16'hbfa7;
mem_array[35087] = 16'h2bfc;
mem_array[35086] = 16'hbf04;
mem_array[35089] = 16'h6314;
mem_array[35088] = 16'hbebb;
mem_array[35091] = 16'h5bef;
mem_array[35090] = 16'hba9b;
mem_array[35093] = 16'h8faa;
mem_array[35092] = 16'hbdad;
mem_array[35095] = 16'h049b;
mem_array[35094] = 16'hbeb9;
mem_array[35097] = 16'hd39b;
mem_array[35096] = 16'h3f49;
mem_array[35099] = 16'h84c0;
mem_array[35098] = 16'hbf0f;
mem_array[35101] = 16'hff6d;
mem_array[35100] = 16'h3f84;
mem_array[35103] = 16'ha2ba;
mem_array[35102] = 16'hbe0c;
mem_array[35105] = 16'h868f;
mem_array[35104] = 16'h3f9b;
mem_array[35107] = 16'h0374;
mem_array[35106] = 16'hbe58;
mem_array[35109] = 16'hcc32;
mem_array[35108] = 16'hbe9a;
mem_array[35111] = 16'h4102;
mem_array[35110] = 16'hbf0c;
mem_array[35113] = 16'h6b09;
mem_array[35112] = 16'h3f1e;
mem_array[35115] = 16'hf2b4;
mem_array[35114] = 16'hbd2b;
mem_array[35117] = 16'h33ae;
mem_array[35116] = 16'hbe42;
mem_array[35119] = 16'h9623;
mem_array[35118] = 16'hbeab;
mem_array[35121] = 16'h7c09;
mem_array[35120] = 16'hbaa9;
mem_array[35123] = 16'h119b;
mem_array[35122] = 16'hbca0;
mem_array[35125] = 16'h1bfb;
mem_array[35124] = 16'hbe82;
mem_array[35127] = 16'hcff1;
mem_array[35126] = 16'h3e85;
mem_array[35129] = 16'h1a39;
mem_array[35128] = 16'h3f3c;
mem_array[35131] = 16'h684c;
mem_array[35130] = 16'hbe3e;
mem_array[35133] = 16'hd5fa;
mem_array[35132] = 16'h3efa;
mem_array[35135] = 16'hc164;
mem_array[35134] = 16'hbeaf;
mem_array[35137] = 16'h05f5;
mem_array[35136] = 16'h3f40;
mem_array[35139] = 16'h1655;
mem_array[35138] = 16'h3c64;
mem_array[35141] = 16'h3349;
mem_array[35140] = 16'hbe6e;
mem_array[35143] = 16'h6995;
mem_array[35142] = 16'h3e31;
mem_array[35145] = 16'hdc03;
mem_array[35144] = 16'hbf83;
mem_array[35147] = 16'ha76d;
mem_array[35146] = 16'h3ea1;
mem_array[35149] = 16'hd4ea;
mem_array[35148] = 16'hbee9;
mem_array[35151] = 16'h4752;
mem_array[35150] = 16'hbd9d;
mem_array[35153] = 16'h3bd7;
mem_array[35152] = 16'h3efa;
mem_array[35155] = 16'hc9f8;
mem_array[35154] = 16'hbece;
mem_array[35157] = 16'hd5cc;
mem_array[35156] = 16'h3f0b;
mem_array[35159] = 16'h3d83;
mem_array[35158] = 16'hbe0b;
mem_array[35161] = 16'heb19;
mem_array[35160] = 16'h3f23;
mem_array[35163] = 16'h12ef;
mem_array[35162] = 16'h3cd2;
mem_array[35165] = 16'h3e4f;
mem_array[35164] = 16'h3fe9;
mem_array[35167] = 16'hb657;
mem_array[35166] = 16'h3f17;
mem_array[35169] = 16'he91f;
mem_array[35168] = 16'hbdf1;
mem_array[35171] = 16'h137f;
mem_array[35170] = 16'h3e1e;
mem_array[35173] = 16'h63d5;
mem_array[35172] = 16'h3f19;
mem_array[35175] = 16'hecf0;
mem_array[35174] = 16'hbd5d;
mem_array[35177] = 16'h2a98;
mem_array[35176] = 16'h3ffc;
mem_array[35179] = 16'hb2e1;
mem_array[35178] = 16'hbc6e;
mem_array[35181] = 16'h4a25;
mem_array[35180] = 16'hbdbf;
mem_array[35183] = 16'hdf8a;
mem_array[35182] = 16'h3d73;
mem_array[35185] = 16'ha5fa;
mem_array[35184] = 16'h3f02;
mem_array[35187] = 16'h9d18;
mem_array[35186] = 16'h3fb7;
mem_array[35189] = 16'h6625;
mem_array[35188] = 16'h3ebb;
mem_array[35191] = 16'h0720;
mem_array[35190] = 16'hbeaf;
mem_array[35193] = 16'h8e0e;
mem_array[35192] = 16'h3f90;
mem_array[35195] = 16'hf729;
mem_array[35194] = 16'h3da6;
mem_array[35197] = 16'h49bc;
mem_array[35196] = 16'hbf35;
mem_array[35199] = 16'h3589;
mem_array[35198] = 16'hbf30;
mem_array[35201] = 16'h49f1;
mem_array[35200] = 16'hbe6a;
mem_array[35203] = 16'h71ec;
mem_array[35202] = 16'hbeae;
mem_array[35205] = 16'h8490;
mem_array[35204] = 16'hbf2b;
mem_array[35207] = 16'h997d;
mem_array[35206] = 16'hbf60;
mem_array[35209] = 16'h47fa;
mem_array[35208] = 16'h3fa0;
mem_array[35211] = 16'hf01e;
mem_array[35210] = 16'h3e81;
mem_array[35213] = 16'h1ad8;
mem_array[35212] = 16'h3ec4;
mem_array[35215] = 16'h1503;
mem_array[35214] = 16'hbd3e;
mem_array[35217] = 16'h10d7;
mem_array[35216] = 16'h3f3f;
mem_array[35219] = 16'ha68d;
mem_array[35218] = 16'hbf15;
mem_array[35221] = 16'h583e;
mem_array[35220] = 16'h3c4e;
mem_array[35223] = 16'h8f28;
mem_array[35222] = 16'hbcf7;
mem_array[35225] = 16'hafea;
mem_array[35224] = 16'h3cc1;
mem_array[35227] = 16'h79f9;
mem_array[35226] = 16'h3cc2;
mem_array[35229] = 16'ha893;
mem_array[35228] = 16'h3b83;
mem_array[35231] = 16'h962d;
mem_array[35230] = 16'hbb35;
mem_array[35233] = 16'h3574;
mem_array[35232] = 16'h3c8a;
mem_array[35235] = 16'heb27;
mem_array[35234] = 16'h3c80;
mem_array[35237] = 16'h48cd;
mem_array[35236] = 16'h3d47;
mem_array[35239] = 16'h58f5;
mem_array[35238] = 16'h3bf3;
mem_array[35241] = 16'hf37a;
mem_array[35240] = 16'hbd1f;
mem_array[35243] = 16'h1232;
mem_array[35242] = 16'h3de8;
mem_array[35245] = 16'hf8b2;
mem_array[35244] = 16'hbd0e;
mem_array[35247] = 16'h1980;
mem_array[35246] = 16'h3d44;
mem_array[35249] = 16'h9928;
mem_array[35248] = 16'h3c9f;
mem_array[35251] = 16'hcc06;
mem_array[35250] = 16'h3bd4;
mem_array[35253] = 16'h0186;
mem_array[35252] = 16'hbbc7;
mem_array[35255] = 16'hf816;
mem_array[35254] = 16'hba30;
mem_array[35257] = 16'h0ecf;
mem_array[35256] = 16'hbd2f;
mem_array[35259] = 16'hf157;
mem_array[35258] = 16'h3cfb;
mem_array[35261] = 16'h1c8c;
mem_array[35260] = 16'hbe0f;
mem_array[35263] = 16'h3379;
mem_array[35262] = 16'h3e65;
mem_array[35265] = 16'h937e;
mem_array[35264] = 16'hbd76;
mem_array[35267] = 16'h26f7;
mem_array[35266] = 16'hbd2b;
mem_array[35269] = 16'h60aa;
mem_array[35268] = 16'hbc8b;
mem_array[35271] = 16'hb14c;
mem_array[35270] = 16'h3cf9;
mem_array[35273] = 16'hc7f7;
mem_array[35272] = 16'h3ea8;
mem_array[35275] = 16'hf25a;
mem_array[35274] = 16'h3e09;
mem_array[35277] = 16'h7ab0;
mem_array[35276] = 16'hbc0a;
mem_array[35279] = 16'hc0cd;
mem_array[35278] = 16'h3dc9;
mem_array[35281] = 16'h6b38;
mem_array[35280] = 16'hbd56;
mem_array[35283] = 16'ha6eb;
mem_array[35282] = 16'h3d64;
mem_array[35285] = 16'hf513;
mem_array[35284] = 16'hbd84;
mem_array[35287] = 16'h6926;
mem_array[35286] = 16'hbd8d;
mem_array[35289] = 16'hf99c;
mem_array[35288] = 16'hbd94;
mem_array[35291] = 16'hf63c;
mem_array[35290] = 16'hbd58;
mem_array[35293] = 16'hd609;
mem_array[35292] = 16'h3c46;
mem_array[35295] = 16'h9260;
mem_array[35294] = 16'h3dbf;
mem_array[35297] = 16'hf0e6;
mem_array[35296] = 16'h3caa;
mem_array[35299] = 16'h8f17;
mem_array[35298] = 16'h3d81;
mem_array[35301] = 16'h2ade;
mem_array[35300] = 16'hbd9a;
mem_array[35303] = 16'h3c60;
mem_array[35302] = 16'hbd5a;
mem_array[35305] = 16'h98ae;
mem_array[35304] = 16'h3d88;
mem_array[35307] = 16'hd0a2;
mem_array[35306] = 16'h3cbd;
mem_array[35309] = 16'h48c4;
mem_array[35308] = 16'h3d11;
mem_array[35311] = 16'hb5c3;
mem_array[35310] = 16'h3df2;
mem_array[35313] = 16'h24df;
mem_array[35312] = 16'hbb45;
mem_array[35315] = 16'h3050;
mem_array[35314] = 16'hbd0a;
mem_array[35317] = 16'h2fc5;
mem_array[35316] = 16'hbd01;
mem_array[35319] = 16'h0373;
mem_array[35318] = 16'hbce3;
mem_array[35321] = 16'h7d8d;
mem_array[35320] = 16'hbd47;
mem_array[35323] = 16'ha230;
mem_array[35322] = 16'h3d81;
mem_array[35325] = 16'h4790;
mem_array[35324] = 16'hbd17;
mem_array[35327] = 16'h783a;
mem_array[35326] = 16'hbb62;
mem_array[35329] = 16'hd0d9;
mem_array[35328] = 16'hbabf;
mem_array[35331] = 16'h6c2d;
mem_array[35330] = 16'h3c4b;
mem_array[35333] = 16'h6442;
mem_array[35332] = 16'h3e0f;
mem_array[35335] = 16'hf445;
mem_array[35334] = 16'hbd8e;
mem_array[35337] = 16'hdafe;
mem_array[35336] = 16'h3d61;
mem_array[35339] = 16'h4754;
mem_array[35338] = 16'h3d2d;
mem_array[35341] = 16'hb664;
mem_array[35340] = 16'hbdd5;
mem_array[35343] = 16'he7d0;
mem_array[35342] = 16'h3d89;
mem_array[35345] = 16'hc1a7;
mem_array[35344] = 16'h3e22;
mem_array[35347] = 16'hdba9;
mem_array[35346] = 16'hbdcf;
mem_array[35349] = 16'h8ed8;
mem_array[35348] = 16'h3cbc;
mem_array[35351] = 16'hdc33;
mem_array[35350] = 16'hbe82;
mem_array[35353] = 16'h6752;
mem_array[35352] = 16'h3e92;
mem_array[35355] = 16'hf0d9;
mem_array[35354] = 16'h3e41;
mem_array[35357] = 16'h83c8;
mem_array[35356] = 16'h3d37;
mem_array[35359] = 16'h5767;
mem_array[35358] = 16'h3d4c;
mem_array[35361] = 16'h3245;
mem_array[35360] = 16'h3c1a;
mem_array[35363] = 16'h5c00;
mem_array[35362] = 16'hbabe;
mem_array[35365] = 16'hbcf7;
mem_array[35364] = 16'hbeb8;
mem_array[35367] = 16'h198c;
mem_array[35366] = 16'h3e8a;
mem_array[35369] = 16'hfd07;
mem_array[35368] = 16'h3eb6;
mem_array[35371] = 16'h2b6e;
mem_array[35370] = 16'h3ecd;
mem_array[35373] = 16'hea1b;
mem_array[35372] = 16'hbcca;
mem_array[35375] = 16'h5979;
mem_array[35374] = 16'h3d0f;
mem_array[35377] = 16'hd97f;
mem_array[35376] = 16'h3d68;
mem_array[35379] = 16'h8098;
mem_array[35378] = 16'h3b88;
mem_array[35381] = 16'h6ffb;
mem_array[35380] = 16'h3e14;
mem_array[35383] = 16'hb231;
mem_array[35382] = 16'h3f0d;
mem_array[35385] = 16'hd805;
mem_array[35384] = 16'h3d43;
mem_array[35387] = 16'h3e58;
mem_array[35386] = 16'hbe23;
mem_array[35389] = 16'h20e3;
mem_array[35388] = 16'h3ec9;
mem_array[35391] = 16'h105f;
mem_array[35390] = 16'hbc2a;
mem_array[35393] = 16'hc942;
mem_array[35392] = 16'h3e30;
mem_array[35395] = 16'h5158;
mem_array[35394] = 16'h3cf9;
mem_array[35397] = 16'h65eb;
mem_array[35396] = 16'hbd86;
mem_array[35399] = 16'ha654;
mem_array[35398] = 16'h3d4d;
mem_array[35401] = 16'h4378;
mem_array[35400] = 16'hbe21;
mem_array[35403] = 16'h6bc1;
mem_array[35402] = 16'h3e32;
mem_array[35405] = 16'h740c;
mem_array[35404] = 16'h3e5c;
mem_array[35407] = 16'h9b4d;
mem_array[35406] = 16'hbe95;
mem_array[35409] = 16'h7b4e;
mem_array[35408] = 16'hbd3d;
mem_array[35411] = 16'h730d;
mem_array[35410] = 16'hbf17;
mem_array[35413] = 16'h25b0;
mem_array[35412] = 16'h3e19;
mem_array[35415] = 16'h4589;
mem_array[35414] = 16'h3e36;
mem_array[35417] = 16'h1a84;
mem_array[35416] = 16'h3f01;
mem_array[35419] = 16'he08e;
mem_array[35418] = 16'hbdc8;
mem_array[35421] = 16'hb366;
mem_array[35420] = 16'hbcc8;
mem_array[35423] = 16'h1355;
mem_array[35422] = 16'hbd13;
mem_array[35425] = 16'h87d5;
mem_array[35424] = 16'hbf44;
mem_array[35427] = 16'h38b6;
mem_array[35426] = 16'h3f5f;
mem_array[35429] = 16'h1be3;
mem_array[35428] = 16'h3d97;
mem_array[35431] = 16'h0559;
mem_array[35430] = 16'h3dbe;
mem_array[35433] = 16'hdd50;
mem_array[35432] = 16'h3ede;
mem_array[35435] = 16'h8f10;
mem_array[35434] = 16'h3ef6;
mem_array[35437] = 16'h072e;
mem_array[35436] = 16'h3d64;
mem_array[35439] = 16'h12d3;
mem_array[35438] = 16'h3df0;
mem_array[35441] = 16'hfce6;
mem_array[35440] = 16'h3dae;
mem_array[35443] = 16'h516b;
mem_array[35442] = 16'h3f42;
mem_array[35445] = 16'h14a0;
mem_array[35444] = 16'h3dc3;
mem_array[35447] = 16'h002f;
mem_array[35446] = 16'h3d25;
mem_array[35449] = 16'hf582;
mem_array[35448] = 16'hbdd3;
mem_array[35451] = 16'h442f;
mem_array[35450] = 16'h3c39;
mem_array[35453] = 16'h0f9e;
mem_array[35452] = 16'hbf22;
mem_array[35455] = 16'hc643;
mem_array[35454] = 16'h3e74;
mem_array[35457] = 16'h8e53;
mem_array[35456] = 16'hbdc3;
mem_array[35459] = 16'h4625;
mem_array[35458] = 16'hbdcf;
mem_array[35461] = 16'h7e97;
mem_array[35460] = 16'hbd70;
mem_array[35463] = 16'hae98;
mem_array[35462] = 16'hbf94;
mem_array[35465] = 16'h2d49;
mem_array[35464] = 16'hbf81;
mem_array[35467] = 16'h3316;
mem_array[35466] = 16'hbf22;
mem_array[35469] = 16'hc2be;
mem_array[35468] = 16'h3f03;
mem_array[35471] = 16'h1280;
mem_array[35470] = 16'hbe93;
mem_array[35473] = 16'hbd09;
mem_array[35472] = 16'hbd54;
mem_array[35475] = 16'hffac;
mem_array[35474] = 16'h3d79;
mem_array[35477] = 16'h3ffe;
mem_array[35476] = 16'h3f29;
mem_array[35479] = 16'h9f80;
mem_array[35478] = 16'h3d4c;
mem_array[35481] = 16'h529d;
mem_array[35480] = 16'hbca1;
mem_array[35483] = 16'hb46c;
mem_array[35482] = 16'h3c0d;
mem_array[35485] = 16'h03bf;
mem_array[35484] = 16'h3e42;
mem_array[35487] = 16'h1078;
mem_array[35486] = 16'h3f34;
mem_array[35489] = 16'h74e9;
mem_array[35488] = 16'h3db3;
mem_array[35491] = 16'he83b;
mem_array[35490] = 16'hbee9;
mem_array[35493] = 16'h16ea;
mem_array[35492] = 16'h3f81;
mem_array[35495] = 16'h6554;
mem_array[35494] = 16'h3d8c;
mem_array[35497] = 16'h2515;
mem_array[35496] = 16'hbf56;
mem_array[35499] = 16'hc902;
mem_array[35498] = 16'hbfa8;
mem_array[35501] = 16'h3cdd;
mem_array[35500] = 16'hbe6a;
mem_array[35503] = 16'hca3e;
mem_array[35502] = 16'h3dd1;
mem_array[35505] = 16'h6f3b;
mem_array[35504] = 16'hbe28;
mem_array[35507] = 16'hfd44;
mem_array[35506] = 16'hbe95;
mem_array[35509] = 16'h4e01;
mem_array[35508] = 16'h3f06;
mem_array[35511] = 16'h6f31;
mem_array[35510] = 16'hbf11;
mem_array[35513] = 16'hf947;
mem_array[35512] = 16'h3dea;
mem_array[35515] = 16'hc823;
mem_array[35514] = 16'hbe91;
mem_array[35517] = 16'h5118;
mem_array[35516] = 16'hbe6b;
mem_array[35519] = 16'h8034;
mem_array[35518] = 16'hbe90;
mem_array[35521] = 16'hbda4;
mem_array[35520] = 16'h3f11;
mem_array[35523] = 16'h5280;
mem_array[35522] = 16'hbef6;
mem_array[35525] = 16'h5894;
mem_array[35524] = 16'hbf18;
mem_array[35527] = 16'h58ad;
mem_array[35526] = 16'h3eb1;
mem_array[35529] = 16'h9448;
mem_array[35528] = 16'h3d8a;
mem_array[35531] = 16'h599b;
mem_array[35530] = 16'h3ec2;
mem_array[35533] = 16'h83d4;
mem_array[35532] = 16'hbd83;
mem_array[35535] = 16'h6d1e;
mem_array[35534] = 16'hbe2a;
mem_array[35537] = 16'ha922;
mem_array[35536] = 16'h3e73;
mem_array[35539] = 16'hda00;
mem_array[35538] = 16'hbf88;
mem_array[35541] = 16'hc0e2;
mem_array[35540] = 16'h3d48;
mem_array[35543] = 16'h9e8f;
mem_array[35542] = 16'hbd50;
mem_array[35545] = 16'hd721;
mem_array[35544] = 16'hbdee;
mem_array[35547] = 16'hbdb0;
mem_array[35546] = 16'hbf10;
mem_array[35549] = 16'h9c32;
mem_array[35548] = 16'hbda8;
mem_array[35551] = 16'h6653;
mem_array[35550] = 16'h3da6;
mem_array[35553] = 16'h8ea0;
mem_array[35552] = 16'hbe9d;
mem_array[35555] = 16'h3692;
mem_array[35554] = 16'hbe5b;
mem_array[35557] = 16'hc04a;
mem_array[35556] = 16'hbfa9;
mem_array[35559] = 16'hc971;
mem_array[35558] = 16'h3e5d;
mem_array[35561] = 16'hbd7d;
mem_array[35560] = 16'h3ed4;
mem_array[35563] = 16'h847a;
mem_array[35562] = 16'h3e0b;
mem_array[35565] = 16'h1daf;
mem_array[35564] = 16'hbee0;
mem_array[35567] = 16'hb500;
mem_array[35566] = 16'h3e8f;
mem_array[35569] = 16'h4531;
mem_array[35568] = 16'h3dad;
mem_array[35571] = 16'h7b52;
mem_array[35570] = 16'hbe5d;
mem_array[35573] = 16'h64cf;
mem_array[35572] = 16'h3e2d;
mem_array[35575] = 16'h26b5;
mem_array[35574] = 16'h3ca1;
mem_array[35577] = 16'h10a8;
mem_array[35576] = 16'hbebf;
mem_array[35579] = 16'hb3ed;
mem_array[35578] = 16'hbf5b;
mem_array[35581] = 16'h1e2a;
mem_array[35580] = 16'hbe27;
mem_array[35583] = 16'hadbb;
mem_array[35582] = 16'hbe19;
mem_array[35585] = 16'hf1c4;
mem_array[35584] = 16'hbd92;
mem_array[35587] = 16'h6e21;
mem_array[35586] = 16'h3d11;
mem_array[35589] = 16'h2fe1;
mem_array[35588] = 16'h3dc4;
mem_array[35591] = 16'hd696;
mem_array[35590] = 16'h3ed3;
mem_array[35593] = 16'hbeff;
mem_array[35592] = 16'hbe11;
mem_array[35595] = 16'heac3;
mem_array[35594] = 16'hbebd;
mem_array[35597] = 16'h670f;
mem_array[35596] = 16'h3d5c;
mem_array[35599] = 16'hc155;
mem_array[35598] = 16'hbf37;
mem_array[35601] = 16'hd58d;
mem_array[35600] = 16'hbdcc;
mem_array[35603] = 16'h742a;
mem_array[35602] = 16'hbcf2;
mem_array[35605] = 16'h0fa1;
mem_array[35604] = 16'h3ee6;
mem_array[35607] = 16'hd7ee;
mem_array[35606] = 16'hbd8a;
mem_array[35609] = 16'ha822;
mem_array[35608] = 16'h3d96;
mem_array[35611] = 16'hbfbe;
mem_array[35610] = 16'h3d07;
mem_array[35613] = 16'h48db;
mem_array[35612] = 16'h3d9e;
mem_array[35615] = 16'hf77a;
mem_array[35614] = 16'h3e60;
mem_array[35617] = 16'hb968;
mem_array[35616] = 16'hbf79;
mem_array[35619] = 16'h1a30;
mem_array[35618] = 16'hbf40;
mem_array[35621] = 16'h33fe;
mem_array[35620] = 16'hbf99;
mem_array[35623] = 16'hab49;
mem_array[35622] = 16'h3d06;
mem_array[35625] = 16'h16fc;
mem_array[35624] = 16'hbed1;
mem_array[35627] = 16'h4e50;
mem_array[35626] = 16'h3cb4;
mem_array[35629] = 16'h75d9;
mem_array[35628] = 16'h3e79;
mem_array[35631] = 16'h6599;
mem_array[35630] = 16'hbf07;
mem_array[35633] = 16'h58cf;
mem_array[35632] = 16'hbe6d;
mem_array[35635] = 16'h7a80;
mem_array[35634] = 16'h3e8e;
mem_array[35637] = 16'hb5f2;
mem_array[35636] = 16'h3c5d;
mem_array[35639] = 16'h1a8d;
mem_array[35638] = 16'hbf3c;
mem_array[35641] = 16'hd832;
mem_array[35640] = 16'hbe69;
mem_array[35643] = 16'hb15f;
mem_array[35642] = 16'hbf75;
mem_array[35645] = 16'h7646;
mem_array[35644] = 16'hbec1;
mem_array[35647] = 16'h8e57;
mem_array[35646] = 16'hbccb;
mem_array[35649] = 16'h9434;
mem_array[35648] = 16'hbe44;
mem_array[35651] = 16'h8cb3;
mem_array[35650] = 16'h3eab;
mem_array[35653] = 16'hd579;
mem_array[35652] = 16'h3e76;
mem_array[35655] = 16'hfd56;
mem_array[35654] = 16'h3dcc;
mem_array[35657] = 16'h2350;
mem_array[35656] = 16'hbe02;
mem_array[35659] = 16'hba39;
mem_array[35658] = 16'hbf32;
mem_array[35661] = 16'hc685;
mem_array[35660] = 16'hbdf9;
mem_array[35663] = 16'hda36;
mem_array[35662] = 16'hbd22;
mem_array[35665] = 16'h90fb;
mem_array[35664] = 16'h3d48;
mem_array[35667] = 16'h28ef;
mem_array[35666] = 16'hbe81;
mem_array[35669] = 16'hac4e;
mem_array[35668] = 16'h3d2e;
mem_array[35671] = 16'h5960;
mem_array[35670] = 16'h3e3c;
mem_array[35673] = 16'hfde1;
mem_array[35672] = 16'h3b5e;
mem_array[35675] = 16'h8d6e;
mem_array[35674] = 16'hbd70;
mem_array[35677] = 16'h1ca4;
mem_array[35676] = 16'hbf21;
mem_array[35679] = 16'hc0d6;
mem_array[35678] = 16'hbf68;
mem_array[35681] = 16'hed74;
mem_array[35680] = 16'hc016;
mem_array[35683] = 16'h409a;
mem_array[35682] = 16'h3e81;
mem_array[35685] = 16'h10e5;
mem_array[35684] = 16'hbeaf;
mem_array[35687] = 16'h67ad;
mem_array[35686] = 16'hbe31;
mem_array[35689] = 16'hbc6f;
mem_array[35688] = 16'h3f0f;
mem_array[35691] = 16'h7dbf;
mem_array[35690] = 16'hbbd6;
mem_array[35693] = 16'h896c;
mem_array[35692] = 16'h3e1a;
mem_array[35695] = 16'hf877;
mem_array[35694] = 16'h3ed4;
mem_array[35697] = 16'h9c66;
mem_array[35696] = 16'h3d0f;
mem_array[35699] = 16'h0a84;
mem_array[35698] = 16'hbf10;
mem_array[35701] = 16'h4416;
mem_array[35700] = 16'hba85;
mem_array[35703] = 16'h64c4;
mem_array[35702] = 16'hbfd4;
mem_array[35705] = 16'haa08;
mem_array[35704] = 16'hbd97;
mem_array[35707] = 16'hf733;
mem_array[35706] = 16'h3c89;
mem_array[35709] = 16'hca9e;
mem_array[35708] = 16'hbe95;
mem_array[35711] = 16'h9e48;
mem_array[35710] = 16'hbdaa;
mem_array[35713] = 16'h95e8;
mem_array[35712] = 16'h3dac;
mem_array[35715] = 16'h8c1b;
mem_array[35714] = 16'h3be6;
mem_array[35717] = 16'h227e;
mem_array[35716] = 16'hbe67;
mem_array[35719] = 16'h9ce5;
mem_array[35718] = 16'h3f07;
mem_array[35721] = 16'h5cbb;
mem_array[35720] = 16'h3cc0;
mem_array[35723] = 16'hb550;
mem_array[35722] = 16'hbd9b;
mem_array[35725] = 16'h71c2;
mem_array[35724] = 16'hbe64;
mem_array[35727] = 16'h8fbf;
mem_array[35726] = 16'hbe69;
mem_array[35729] = 16'h242d;
mem_array[35728] = 16'hbde4;
mem_array[35731] = 16'h3211;
mem_array[35730] = 16'hbd4f;
mem_array[35733] = 16'h584b;
mem_array[35732] = 16'h3ee2;
mem_array[35735] = 16'h8822;
mem_array[35734] = 16'hbeb8;
mem_array[35737] = 16'h9f3f;
mem_array[35736] = 16'hbf2c;
mem_array[35739] = 16'h3ccc;
mem_array[35738] = 16'hbe6b;
mem_array[35741] = 16'h02f3;
mem_array[35740] = 16'hbe3a;
mem_array[35743] = 16'hbb08;
mem_array[35742] = 16'h3dec;
mem_array[35745] = 16'h731d;
mem_array[35744] = 16'hbe43;
mem_array[35747] = 16'h571a;
mem_array[35746] = 16'hbe21;
mem_array[35749] = 16'he476;
mem_array[35748] = 16'h3dcc;
mem_array[35751] = 16'ha4be;
mem_array[35750] = 16'hbf23;
mem_array[35753] = 16'h938b;
mem_array[35752] = 16'h3e36;
mem_array[35755] = 16'h3b7b;
mem_array[35754] = 16'h3d92;
mem_array[35757] = 16'h8094;
mem_array[35756] = 16'hbe63;
mem_array[35759] = 16'h7aab;
mem_array[35758] = 16'hbeb7;
mem_array[35761] = 16'h457b;
mem_array[35760] = 16'hbe28;
mem_array[35763] = 16'h914a;
mem_array[35762] = 16'hbf7b;
mem_array[35765] = 16'h7ba8;
mem_array[35764] = 16'hbdbe;
mem_array[35767] = 16'h21ec;
mem_array[35766] = 16'hbd31;
mem_array[35769] = 16'h594d;
mem_array[35768] = 16'h3e4e;
mem_array[35771] = 16'h2dbb;
mem_array[35770] = 16'hbd25;
mem_array[35773] = 16'hb93e;
mem_array[35772] = 16'hbd06;
mem_array[35775] = 16'h9650;
mem_array[35774] = 16'hbe06;
mem_array[35777] = 16'h3aae;
mem_array[35776] = 16'hbcd4;
mem_array[35779] = 16'h884d;
mem_array[35778] = 16'hbe5c;
mem_array[35781] = 16'hb7dc;
mem_array[35780] = 16'hbda7;
mem_array[35783] = 16'h3bf4;
mem_array[35782] = 16'hbd4e;
mem_array[35785] = 16'hc8cd;
mem_array[35784] = 16'hbeee;
mem_array[35787] = 16'hf605;
mem_array[35786] = 16'hbdde;
mem_array[35789] = 16'h9790;
mem_array[35788] = 16'h3e16;
mem_array[35791] = 16'h23b3;
mem_array[35790] = 16'hbd88;
mem_array[35793] = 16'h82d9;
mem_array[35792] = 16'hbe9d;
mem_array[35795] = 16'h7736;
mem_array[35794] = 16'hbe7f;
mem_array[35797] = 16'ha716;
mem_array[35796] = 16'hbf80;
mem_array[35799] = 16'h1faa;
mem_array[35798] = 16'hbe95;
mem_array[35801] = 16'hcf6b;
mem_array[35800] = 16'h3f55;
mem_array[35803] = 16'he057;
mem_array[35802] = 16'h3e37;
mem_array[35805] = 16'h01ba;
mem_array[35804] = 16'hbdd7;
mem_array[35807] = 16'hb057;
mem_array[35806] = 16'hbdb9;
mem_array[35809] = 16'h41b8;
mem_array[35808] = 16'hbd41;
mem_array[35811] = 16'hf4fe;
mem_array[35810] = 16'hbf2f;
mem_array[35813] = 16'h415d;
mem_array[35812] = 16'h3df1;
mem_array[35815] = 16'hab36;
mem_array[35814] = 16'h3d4e;
mem_array[35817] = 16'h8736;
mem_array[35816] = 16'hbe49;
mem_array[35819] = 16'hd767;
mem_array[35818] = 16'h3de2;
mem_array[35821] = 16'h7728;
mem_array[35820] = 16'hbdce;
mem_array[35823] = 16'h89e6;
mem_array[35822] = 16'h3e10;
mem_array[35825] = 16'h4dfb;
mem_array[35824] = 16'hbd37;
mem_array[35827] = 16'h812f;
mem_array[35826] = 16'h3dc3;
mem_array[35829] = 16'h6bb4;
mem_array[35828] = 16'h3f00;
mem_array[35831] = 16'hc1d6;
mem_array[35830] = 16'h3de3;
mem_array[35833] = 16'hfbc5;
mem_array[35832] = 16'hbd92;
mem_array[35835] = 16'h25c3;
mem_array[35834] = 16'hbd79;
mem_array[35837] = 16'h0f03;
mem_array[35836] = 16'h3dcc;
mem_array[35839] = 16'h19a3;
mem_array[35838] = 16'h3e85;
mem_array[35841] = 16'hc58c;
mem_array[35840] = 16'hbd67;
mem_array[35843] = 16'h2e9f;
mem_array[35842] = 16'hbd32;
mem_array[35845] = 16'h9307;
mem_array[35844] = 16'hbe50;
mem_array[35847] = 16'h7ddf;
mem_array[35846] = 16'h3d90;
mem_array[35849] = 16'h661e;
mem_array[35848] = 16'h3e70;
mem_array[35851] = 16'hbafe;
mem_array[35850] = 16'hbe1a;
mem_array[35853] = 16'h9101;
mem_array[35852] = 16'h3e1b;
mem_array[35855] = 16'ha8db;
mem_array[35854] = 16'hbe77;
mem_array[35857] = 16'hfbf9;
mem_array[35856] = 16'hbf68;
mem_array[35859] = 16'h2053;
mem_array[35858] = 16'hbfa1;
mem_array[35861] = 16'h1a13;
mem_array[35860] = 16'h3f14;
mem_array[35863] = 16'h63e9;
mem_array[35862] = 16'h3e18;
mem_array[35865] = 16'hac13;
mem_array[35864] = 16'hbd80;
mem_array[35867] = 16'hc22c;
mem_array[35866] = 16'hbde6;
mem_array[35869] = 16'he383;
mem_array[35868] = 16'hbd58;
mem_array[35871] = 16'he14c;
mem_array[35870] = 16'hbe8d;
mem_array[35873] = 16'hc070;
mem_array[35872] = 16'h3dfb;
mem_array[35875] = 16'h994b;
mem_array[35874] = 16'h3aad;
mem_array[35877] = 16'haf1c;
mem_array[35876] = 16'hbbc2;
mem_array[35879] = 16'hb97a;
mem_array[35878] = 16'hbe08;
mem_array[35881] = 16'h8806;
mem_array[35880] = 16'h3d96;
mem_array[35883] = 16'hf40b;
mem_array[35882] = 16'hbdf3;
mem_array[35885] = 16'h4096;
mem_array[35884] = 16'h3e00;
mem_array[35887] = 16'h83e3;
mem_array[35886] = 16'h3e8b;
mem_array[35889] = 16'h8b73;
mem_array[35888] = 16'h3e58;
mem_array[35891] = 16'ha0da;
mem_array[35890] = 16'h3d7d;
mem_array[35893] = 16'h7bbd;
mem_array[35892] = 16'hbd35;
mem_array[35895] = 16'hbf6c;
mem_array[35894] = 16'hbd9b;
mem_array[35897] = 16'hf2fa;
mem_array[35896] = 16'h3dd3;
mem_array[35899] = 16'hbf07;
mem_array[35898] = 16'h3e4c;
mem_array[35901] = 16'hcec3;
mem_array[35900] = 16'hbd6a;
mem_array[35903] = 16'hfc1d;
mem_array[35902] = 16'hbb3a;
mem_array[35905] = 16'hcfaf;
mem_array[35904] = 16'h3ddf;
mem_array[35907] = 16'hd00c;
mem_array[35906] = 16'hbc9e;
mem_array[35909] = 16'h3724;
mem_array[35908] = 16'h3e4c;
mem_array[35911] = 16'h7871;
mem_array[35910] = 16'hbd70;
mem_array[35913] = 16'h3994;
mem_array[35912] = 16'hbb95;
mem_array[35915] = 16'hcca4;
mem_array[35914] = 16'hbe69;
mem_array[35917] = 16'hd380;
mem_array[35916] = 16'hbf23;
mem_array[35919] = 16'h9e23;
mem_array[35918] = 16'hbf8f;
mem_array[35921] = 16'hf7ea;
mem_array[35920] = 16'h3e8a;
mem_array[35923] = 16'hae11;
mem_array[35922] = 16'hbb6f;
mem_array[35925] = 16'he024;
mem_array[35924] = 16'hbdd1;
mem_array[35927] = 16'h4097;
mem_array[35926] = 16'hbecc;
mem_array[35929] = 16'h0635;
mem_array[35928] = 16'h3e81;
mem_array[35931] = 16'hfd68;
mem_array[35930] = 16'h3e1c;
mem_array[35933] = 16'h8e4a;
mem_array[35932] = 16'h3e0a;
mem_array[35935] = 16'h6c8e;
mem_array[35934] = 16'hbc76;
mem_array[35937] = 16'h1932;
mem_array[35936] = 16'h3e3b;
mem_array[35939] = 16'hc17d;
mem_array[35938] = 16'h3da3;
mem_array[35941] = 16'h5124;
mem_array[35940] = 16'hbe55;
mem_array[35943] = 16'ha9cd;
mem_array[35942] = 16'h3d59;
mem_array[35945] = 16'hf288;
mem_array[35944] = 16'h3cf9;
mem_array[35947] = 16'he932;
mem_array[35946] = 16'h3ecb;
mem_array[35949] = 16'ha529;
mem_array[35948] = 16'h3c53;
mem_array[35951] = 16'hc19b;
mem_array[35950] = 16'h3d8c;
mem_array[35953] = 16'h5734;
mem_array[35952] = 16'h3dbb;
mem_array[35955] = 16'h6a0d;
mem_array[35954] = 16'hbe2f;
mem_array[35957] = 16'h039a;
mem_array[35956] = 16'hbe39;
mem_array[35959] = 16'h3cf6;
mem_array[35958] = 16'h3c99;
mem_array[35961] = 16'h73f5;
mem_array[35960] = 16'hbdd7;
mem_array[35963] = 16'h93d3;
mem_array[35962] = 16'h3b97;
mem_array[35965] = 16'h677b;
mem_array[35964] = 16'hbcba;
mem_array[35967] = 16'h5323;
mem_array[35966] = 16'hbd0b;
mem_array[35969] = 16'heb62;
mem_array[35968] = 16'hbee0;
mem_array[35971] = 16'h198c;
mem_array[35970] = 16'hbe29;
mem_array[35973] = 16'h0197;
mem_array[35972] = 16'hbe40;
mem_array[35975] = 16'h7d4e;
mem_array[35974] = 16'hbe01;
mem_array[35977] = 16'hee81;
mem_array[35976] = 16'hbef8;
mem_array[35979] = 16'h790a;
mem_array[35978] = 16'hbf1a;
mem_array[35981] = 16'hb44a;
mem_array[35980] = 16'h3e94;
mem_array[35983] = 16'ha0a8;
mem_array[35982] = 16'h3aab;
mem_array[35985] = 16'h1287;
mem_array[35984] = 16'h3af7;
mem_array[35987] = 16'h3a8b;
mem_array[35986] = 16'hbca2;
mem_array[35989] = 16'h32ca;
mem_array[35988] = 16'hbe79;
mem_array[35991] = 16'h8c51;
mem_array[35990] = 16'hbd9b;
mem_array[35993] = 16'h0848;
mem_array[35992] = 16'hbdc3;
mem_array[35995] = 16'hf45e;
mem_array[35994] = 16'h3e0f;
mem_array[35997] = 16'h46ab;
mem_array[35996] = 16'hbe17;
mem_array[35999] = 16'h2e59;
mem_array[35998] = 16'h3e6e;
mem_array[36001] = 16'h0f3f;
mem_array[36000] = 16'hbca4;
mem_array[36003] = 16'h1a27;
mem_array[36002] = 16'hbd8d;
mem_array[36005] = 16'h994e;
mem_array[36004] = 16'h3dc2;
mem_array[36007] = 16'h45ee;
mem_array[36006] = 16'h3d4e;
mem_array[36009] = 16'h8da2;
mem_array[36008] = 16'hbe85;
mem_array[36011] = 16'hed1d;
mem_array[36010] = 16'hbe00;
mem_array[36013] = 16'h3ba4;
mem_array[36012] = 16'h3e21;
mem_array[36015] = 16'h1571;
mem_array[36014] = 16'hbc0b;
mem_array[36017] = 16'h936d;
mem_array[36016] = 16'h3d74;
mem_array[36019] = 16'ha84b;
mem_array[36018] = 16'h3e32;
mem_array[36021] = 16'h99c9;
mem_array[36020] = 16'hbc1a;
mem_array[36023] = 16'h3ba5;
mem_array[36022] = 16'hbd82;
mem_array[36025] = 16'he4f2;
mem_array[36024] = 16'h3db6;
mem_array[36027] = 16'hf3a7;
mem_array[36026] = 16'hbda1;
mem_array[36029] = 16'h2bad;
mem_array[36028] = 16'hbea4;
mem_array[36031] = 16'hfa54;
mem_array[36030] = 16'hbe7c;
mem_array[36033] = 16'h8315;
mem_array[36032] = 16'hbd10;
mem_array[36035] = 16'hff2c;
mem_array[36034] = 16'h3dca;
mem_array[36037] = 16'h7915;
mem_array[36036] = 16'hbe67;
mem_array[36039] = 16'hb2a1;
mem_array[36038] = 16'hbe1a;
mem_array[36041] = 16'hb08e;
mem_array[36040] = 16'hbdb2;
mem_array[36043] = 16'h265b;
mem_array[36042] = 16'hbdcd;
mem_array[36045] = 16'hef76;
mem_array[36044] = 16'h3e51;
mem_array[36047] = 16'h3e7c;
mem_array[36046] = 16'hbea3;
mem_array[36049] = 16'h56b0;
mem_array[36048] = 16'hbbb0;
mem_array[36051] = 16'h0840;
mem_array[36050] = 16'hbeba;
mem_array[36053] = 16'h99ff;
mem_array[36052] = 16'hbe11;
mem_array[36055] = 16'h50f0;
mem_array[36054] = 16'h3d14;
mem_array[36057] = 16'hf052;
mem_array[36056] = 16'hbe8b;
mem_array[36059] = 16'h6b0c;
mem_array[36058] = 16'h3e9b;
mem_array[36061] = 16'h0622;
mem_array[36060] = 16'hbe26;
mem_array[36063] = 16'h7134;
mem_array[36062] = 16'h3e0a;
mem_array[36065] = 16'h5811;
mem_array[36064] = 16'h3b88;
mem_array[36067] = 16'hffb2;
mem_array[36066] = 16'hbe29;
mem_array[36069] = 16'ha547;
mem_array[36068] = 16'hbea4;
mem_array[36071] = 16'h8a82;
mem_array[36070] = 16'h3d69;
mem_array[36073] = 16'h65e6;
mem_array[36072] = 16'h3e1f;
mem_array[36075] = 16'h35d4;
mem_array[36074] = 16'hbd81;
mem_array[36077] = 16'hac99;
mem_array[36076] = 16'hbdef;
mem_array[36079] = 16'h7d3d;
mem_array[36078] = 16'h3e4d;
mem_array[36081] = 16'h9863;
mem_array[36080] = 16'hbc8d;
mem_array[36083] = 16'hfe84;
mem_array[36082] = 16'hbc6a;
mem_array[36085] = 16'h6b44;
mem_array[36084] = 16'hbd8f;
mem_array[36087] = 16'h6d67;
mem_array[36086] = 16'hbec8;
mem_array[36089] = 16'hb55f;
mem_array[36088] = 16'h3dc4;
mem_array[36091] = 16'hd4c7;
mem_array[36090] = 16'hbe01;
mem_array[36093] = 16'hd0f1;
mem_array[36092] = 16'hbe02;
mem_array[36095] = 16'h65a9;
mem_array[36094] = 16'h3d29;
mem_array[36097] = 16'hb3f0;
mem_array[36096] = 16'hbea2;
mem_array[36099] = 16'h6509;
mem_array[36098] = 16'hbd9c;
mem_array[36101] = 16'h7df4;
mem_array[36100] = 16'hbe40;
mem_array[36103] = 16'he94e;
mem_array[36102] = 16'h3ed6;
mem_array[36105] = 16'hf6a8;
mem_array[36104] = 16'h3f03;
mem_array[36107] = 16'hbc25;
mem_array[36106] = 16'hbcce;
mem_array[36109] = 16'h3ba3;
mem_array[36108] = 16'h3df4;
mem_array[36111] = 16'haa3b;
mem_array[36110] = 16'hbe16;
mem_array[36113] = 16'h48b5;
mem_array[36112] = 16'h3d9e;
mem_array[36115] = 16'h6f04;
mem_array[36114] = 16'h3d9d;
mem_array[36117] = 16'h03d0;
mem_array[36116] = 16'hbef0;
mem_array[36119] = 16'hb2ab;
mem_array[36118] = 16'h3e8b;
mem_array[36121] = 16'ha45b;
mem_array[36120] = 16'hbea4;
mem_array[36123] = 16'h064e;
mem_array[36122] = 16'hbd21;
mem_array[36125] = 16'h5409;
mem_array[36124] = 16'h3dc9;
mem_array[36127] = 16'h59f5;
mem_array[36126] = 16'hbbc6;
mem_array[36129] = 16'hb366;
mem_array[36128] = 16'hbfaf;
mem_array[36131] = 16'ha175;
mem_array[36130] = 16'hbca5;
mem_array[36133] = 16'hf9e1;
mem_array[36132] = 16'h3e3d;
mem_array[36135] = 16'h7ce2;
mem_array[36134] = 16'h3d5f;
mem_array[36137] = 16'h0b83;
mem_array[36136] = 16'hbe90;
mem_array[36139] = 16'h9783;
mem_array[36138] = 16'hbdc2;
mem_array[36141] = 16'h8f15;
mem_array[36140] = 16'hbdc7;
mem_array[36143] = 16'hf736;
mem_array[36142] = 16'h3d33;
mem_array[36145] = 16'hec72;
mem_array[36144] = 16'hbb41;
mem_array[36147] = 16'hc8d2;
mem_array[36146] = 16'hbeb7;
mem_array[36149] = 16'h11c6;
mem_array[36148] = 16'h3daf;
mem_array[36151] = 16'h568f;
mem_array[36150] = 16'hbdd6;
mem_array[36153] = 16'h2427;
mem_array[36152] = 16'hbd9a;
mem_array[36155] = 16'hbcfc;
mem_array[36154] = 16'h3d11;
mem_array[36157] = 16'hd148;
mem_array[36156] = 16'hbeb2;
mem_array[36159] = 16'h4e71;
mem_array[36158] = 16'hbdd6;
mem_array[36161] = 16'h2334;
mem_array[36160] = 16'hbe38;
mem_array[36163] = 16'h7a5c;
mem_array[36162] = 16'h3dc3;
mem_array[36165] = 16'h7ee4;
mem_array[36164] = 16'h3e93;
mem_array[36167] = 16'heac5;
mem_array[36166] = 16'h3c24;
mem_array[36169] = 16'h68cb;
mem_array[36168] = 16'hb938;
mem_array[36171] = 16'h9031;
mem_array[36170] = 16'hbcce;
mem_array[36173] = 16'hfffa;
mem_array[36172] = 16'h3d8b;
mem_array[36175] = 16'h43d7;
mem_array[36174] = 16'hbe25;
mem_array[36177] = 16'h74b9;
mem_array[36176] = 16'hbf69;
mem_array[36179] = 16'h4a5c;
mem_array[36178] = 16'h3c3b;
mem_array[36181] = 16'h118a;
mem_array[36180] = 16'hbef7;
mem_array[36183] = 16'hb8cd;
mem_array[36182] = 16'hbea7;
mem_array[36185] = 16'hf883;
mem_array[36184] = 16'hbd8e;
mem_array[36187] = 16'h2876;
mem_array[36186] = 16'h3df3;
mem_array[36189] = 16'h3447;
mem_array[36188] = 16'hbf81;
mem_array[36191] = 16'haad3;
mem_array[36190] = 16'h3c2d;
mem_array[36193] = 16'h04d9;
mem_array[36192] = 16'hbcf0;
mem_array[36195] = 16'hfb2c;
mem_array[36194] = 16'hbd4c;
mem_array[36197] = 16'h8bfb;
mem_array[36196] = 16'hbe92;
mem_array[36199] = 16'hb8f6;
mem_array[36198] = 16'h3e5f;
mem_array[36201] = 16'h2d0f;
mem_array[36200] = 16'hbd6f;
mem_array[36203] = 16'h4cdf;
mem_array[36202] = 16'hbd3e;
mem_array[36205] = 16'h1e6a;
mem_array[36204] = 16'hbd6d;
mem_array[36207] = 16'h321a;
mem_array[36206] = 16'h3c95;
mem_array[36209] = 16'hdb5d;
mem_array[36208] = 16'h3f03;
mem_array[36211] = 16'h0441;
mem_array[36210] = 16'hbd8f;
mem_array[36213] = 16'h83e6;
mem_array[36212] = 16'h3dcd;
mem_array[36215] = 16'h11ab;
mem_array[36214] = 16'h3e8e;
mem_array[36217] = 16'ha7fc;
mem_array[36216] = 16'hbee8;
mem_array[36219] = 16'h3640;
mem_array[36218] = 16'hbc59;
mem_array[36221] = 16'h6486;
mem_array[36220] = 16'hbe59;
mem_array[36223] = 16'h67aa;
mem_array[36222] = 16'h3bf6;
mem_array[36225] = 16'h6765;
mem_array[36224] = 16'h3ce8;
mem_array[36227] = 16'h6c0c;
mem_array[36226] = 16'hbe06;
mem_array[36229] = 16'h2889;
mem_array[36228] = 16'hbd41;
mem_array[36231] = 16'h6bc5;
mem_array[36230] = 16'hbe67;
mem_array[36233] = 16'h76fc;
mem_array[36232] = 16'h3e1f;
mem_array[36235] = 16'hb8f0;
mem_array[36234] = 16'hbc98;
mem_array[36237] = 16'ha075;
mem_array[36236] = 16'hbf3b;
mem_array[36239] = 16'hb36f;
mem_array[36238] = 16'h3e53;
mem_array[36241] = 16'hdda7;
mem_array[36240] = 16'hbf26;
mem_array[36243] = 16'h2837;
mem_array[36242] = 16'h3983;
mem_array[36245] = 16'hd994;
mem_array[36244] = 16'hbca1;
mem_array[36247] = 16'hc1f4;
mem_array[36246] = 16'hbe60;
mem_array[36249] = 16'hd06c;
mem_array[36248] = 16'hbfde;
mem_array[36251] = 16'h7750;
mem_array[36250] = 16'h3e40;
mem_array[36253] = 16'hbf43;
mem_array[36252] = 16'h3dfb;
mem_array[36255] = 16'hc02f;
mem_array[36254] = 16'hbe26;
mem_array[36257] = 16'h36c8;
mem_array[36256] = 16'hbebc;
mem_array[36259] = 16'hd96e;
mem_array[36258] = 16'h3ea3;
mem_array[36261] = 16'h84fd;
mem_array[36260] = 16'h3ae1;
mem_array[36263] = 16'h4664;
mem_array[36262] = 16'h3dbb;
mem_array[36265] = 16'h6879;
mem_array[36264] = 16'hbd0d;
mem_array[36267] = 16'hdb0a;
mem_array[36266] = 16'h3ccc;
mem_array[36269] = 16'h1928;
mem_array[36268] = 16'h3e8d;
mem_array[36271] = 16'h9fed;
mem_array[36270] = 16'hbdcc;
mem_array[36273] = 16'h13b0;
mem_array[36272] = 16'h3d1c;
mem_array[36275] = 16'h6511;
mem_array[36274] = 16'hbe6d;
mem_array[36277] = 16'h12a2;
mem_array[36276] = 16'hbe67;
mem_array[36279] = 16'h4d55;
mem_array[36278] = 16'hbdf1;
mem_array[36281] = 16'h73d9;
mem_array[36280] = 16'hbd1b;
mem_array[36283] = 16'h1590;
mem_array[36282] = 16'hbc0b;
mem_array[36285] = 16'hdad0;
mem_array[36284] = 16'h3e2a;
mem_array[36287] = 16'h577c;
mem_array[36286] = 16'hbc60;
mem_array[36289] = 16'h8e35;
mem_array[36288] = 16'hbe88;
mem_array[36291] = 16'h64b4;
mem_array[36290] = 16'hbd94;
mem_array[36293] = 16'h7004;
mem_array[36292] = 16'h3e3b;
mem_array[36295] = 16'hb9b9;
mem_array[36294] = 16'h3e1c;
mem_array[36297] = 16'h51c5;
mem_array[36296] = 16'hbf6a;
mem_array[36299] = 16'he42b;
mem_array[36298] = 16'h3e2d;
mem_array[36301] = 16'h3dda;
mem_array[36300] = 16'h3dd3;
mem_array[36303] = 16'hb461;
mem_array[36302] = 16'h3e43;
mem_array[36305] = 16'h357c;
mem_array[36304] = 16'h3e60;
mem_array[36307] = 16'hd41e;
mem_array[36306] = 16'hbe22;
mem_array[36309] = 16'hfd60;
mem_array[36308] = 16'hbfd2;
mem_array[36311] = 16'h4cb2;
mem_array[36310] = 16'h3e78;
mem_array[36313] = 16'h5b24;
mem_array[36312] = 16'hbe9c;
mem_array[36315] = 16'h5a27;
mem_array[36314] = 16'hbdd5;
mem_array[36317] = 16'h125b;
mem_array[36316] = 16'hbf1a;
mem_array[36319] = 16'he0e1;
mem_array[36318] = 16'hbefb;
mem_array[36321] = 16'haffb;
mem_array[36320] = 16'hbc88;
mem_array[36323] = 16'he7cb;
mem_array[36322] = 16'hbc95;
mem_array[36325] = 16'h2fd5;
mem_array[36324] = 16'h3d6d;
mem_array[36327] = 16'hece4;
mem_array[36326] = 16'hbe02;
mem_array[36329] = 16'h0a36;
mem_array[36328] = 16'h3eb1;
mem_array[36331] = 16'h49c4;
mem_array[36330] = 16'h3e48;
mem_array[36333] = 16'hb073;
mem_array[36332] = 16'h3dad;
mem_array[36335] = 16'h32a2;
mem_array[36334] = 16'h3e4b;
mem_array[36337] = 16'hb627;
mem_array[36336] = 16'hbec0;
mem_array[36339] = 16'h106d;
mem_array[36338] = 16'h3e7a;
mem_array[36341] = 16'h189e;
mem_array[36340] = 16'hbe7f;
mem_array[36343] = 16'h8c49;
mem_array[36342] = 16'hbd4b;
mem_array[36345] = 16'h9e0a;
mem_array[36344] = 16'hbc99;
mem_array[36347] = 16'h00f4;
mem_array[36346] = 16'hbb8a;
mem_array[36349] = 16'hb9c6;
mem_array[36348] = 16'hbe8f;
mem_array[36351] = 16'hbdc0;
mem_array[36350] = 16'hbe80;
mem_array[36353] = 16'h2661;
mem_array[36352] = 16'h3e13;
mem_array[36355] = 16'he790;
mem_array[36354] = 16'hbdef;
mem_array[36357] = 16'hc898;
mem_array[36356] = 16'hbf48;
mem_array[36359] = 16'hb55a;
mem_array[36358] = 16'h3e33;
mem_array[36361] = 16'h23c6;
mem_array[36360] = 16'hbf33;
mem_array[36363] = 16'h0197;
mem_array[36362] = 16'h3d9f;
mem_array[36365] = 16'h0334;
mem_array[36364] = 16'h3d54;
mem_array[36367] = 16'h759d;
mem_array[36366] = 16'hbea1;
mem_array[36369] = 16'h0482;
mem_array[36368] = 16'hbde7;
mem_array[36371] = 16'h787a;
mem_array[36370] = 16'h3d9d;
mem_array[36373] = 16'h086a;
mem_array[36372] = 16'hbd08;
mem_array[36375] = 16'ha8d4;
mem_array[36374] = 16'hbdee;
mem_array[36377] = 16'hc17a;
mem_array[36376] = 16'h3e1b;
mem_array[36379] = 16'ha13a;
mem_array[36378] = 16'h3e81;
mem_array[36381] = 16'ha914;
mem_array[36380] = 16'hbd70;
mem_array[36383] = 16'hf069;
mem_array[36382] = 16'h3d19;
mem_array[36385] = 16'hc30c;
mem_array[36384] = 16'hbdd8;
mem_array[36387] = 16'hde87;
mem_array[36386] = 16'h3d60;
mem_array[36389] = 16'hecf8;
mem_array[36388] = 16'hbd7b;
mem_array[36391] = 16'h96c9;
mem_array[36390] = 16'h3e1e;
mem_array[36393] = 16'h643d;
mem_array[36392] = 16'h3d99;
mem_array[36395] = 16'h96ca;
mem_array[36394] = 16'hbc74;
mem_array[36397] = 16'hb63b;
mem_array[36396] = 16'hbe93;
mem_array[36399] = 16'h0656;
mem_array[36398] = 16'h3e16;
mem_array[36401] = 16'h3488;
mem_array[36400] = 16'h3e10;
mem_array[36403] = 16'h5927;
mem_array[36402] = 16'h3dc5;
mem_array[36405] = 16'h897b;
mem_array[36404] = 16'hbc64;
mem_array[36407] = 16'h78bb;
mem_array[36406] = 16'hbdcd;
mem_array[36409] = 16'h2f1c;
mem_array[36408] = 16'hbdcb;
mem_array[36411] = 16'had49;
mem_array[36410] = 16'hbf3b;
mem_array[36413] = 16'hafb5;
mem_array[36412] = 16'h3e45;
mem_array[36415] = 16'h69f1;
mem_array[36414] = 16'hbe18;
mem_array[36417] = 16'he4b7;
mem_array[36416] = 16'hbe38;
mem_array[36419] = 16'hde2f;
mem_array[36418] = 16'hbbc4;
mem_array[36421] = 16'h4084;
mem_array[36420] = 16'h3d90;
mem_array[36423] = 16'hc570;
mem_array[36422] = 16'h3d21;
mem_array[36425] = 16'h9a5a;
mem_array[36424] = 16'h3d61;
mem_array[36427] = 16'hfda8;
mem_array[36426] = 16'hbedd;
mem_array[36429] = 16'h8455;
mem_array[36428] = 16'hbe55;
mem_array[36431] = 16'h8921;
mem_array[36430] = 16'hbdf1;
mem_array[36433] = 16'h1db4;
mem_array[36432] = 16'hbda3;
mem_array[36435] = 16'h26a9;
mem_array[36434] = 16'hbddc;
mem_array[36437] = 16'ha7ad;
mem_array[36436] = 16'hbee1;
mem_array[36439] = 16'hb10e;
mem_array[36438] = 16'h3d06;
mem_array[36441] = 16'h8a48;
mem_array[36440] = 16'hbdfc;
mem_array[36443] = 16'h0544;
mem_array[36442] = 16'hbd3a;
mem_array[36445] = 16'h0ba5;
mem_array[36444] = 16'hbf02;
mem_array[36447] = 16'h5c80;
mem_array[36446] = 16'h3ebb;
mem_array[36449] = 16'h22c1;
mem_array[36448] = 16'h3d8a;
mem_array[36451] = 16'hb2ec;
mem_array[36450] = 16'h3cf6;
mem_array[36453] = 16'hde92;
mem_array[36452] = 16'h3ef7;
mem_array[36455] = 16'hf379;
mem_array[36454] = 16'hbdd4;
mem_array[36457] = 16'h2bfc;
mem_array[36456] = 16'hbf1b;
mem_array[36459] = 16'h7f9b;
mem_array[36458] = 16'hbe03;
mem_array[36461] = 16'h50ac;
mem_array[36460] = 16'hbd03;
mem_array[36463] = 16'hb407;
mem_array[36462] = 16'hbdb9;
mem_array[36465] = 16'h47d8;
mem_array[36464] = 16'h3e13;
mem_array[36467] = 16'h0766;
mem_array[36466] = 16'hbd8c;
mem_array[36469] = 16'h3d02;
mem_array[36468] = 16'hbe3c;
mem_array[36471] = 16'h7cb5;
mem_array[36470] = 16'hbf7e;
mem_array[36473] = 16'h584e;
mem_array[36472] = 16'h3e3c;
mem_array[36475] = 16'h31ae;
mem_array[36474] = 16'h3dd4;
mem_array[36477] = 16'ha77e;
mem_array[36476] = 16'h3e48;
mem_array[36479] = 16'h7219;
mem_array[36478] = 16'h3e96;
mem_array[36481] = 16'h997c;
mem_array[36480] = 16'hbf5d;
mem_array[36483] = 16'h2423;
mem_array[36482] = 16'hbe77;
mem_array[36485] = 16'hd258;
mem_array[36484] = 16'hbb91;
mem_array[36487] = 16'hbddc;
mem_array[36486] = 16'hbea7;
mem_array[36489] = 16'hd059;
mem_array[36488] = 16'h3ed9;
mem_array[36491] = 16'h2d13;
mem_array[36490] = 16'hbdd8;
mem_array[36493] = 16'hec69;
mem_array[36492] = 16'hbe32;
mem_array[36495] = 16'h6cb5;
mem_array[36494] = 16'hbe7f;
mem_array[36497] = 16'hf62e;
mem_array[36496] = 16'hbe62;
mem_array[36499] = 16'h5dcc;
mem_array[36498] = 16'h3e7c;
mem_array[36501] = 16'hda93;
mem_array[36500] = 16'h3dfd;
mem_array[36503] = 16'hc4ce;
mem_array[36502] = 16'hbd97;
mem_array[36505] = 16'h2b9c;
mem_array[36504] = 16'hbf18;
mem_array[36507] = 16'h0cad;
mem_array[36506] = 16'h3ec7;
mem_array[36509] = 16'h43c3;
mem_array[36508] = 16'h3e1f;
mem_array[36511] = 16'h0847;
mem_array[36510] = 16'hbd43;
mem_array[36513] = 16'h30f6;
mem_array[36512] = 16'h3e50;
mem_array[36515] = 16'hf33d;
mem_array[36514] = 16'h3f0e;
mem_array[36517] = 16'h50e7;
mem_array[36516] = 16'hbf0f;
mem_array[36519] = 16'he3fa;
mem_array[36518] = 16'h3edc;
mem_array[36521] = 16'h23a1;
mem_array[36520] = 16'hbe3d;
mem_array[36523] = 16'hbe19;
mem_array[36522] = 16'h3df5;
mem_array[36525] = 16'ha8fb;
mem_array[36524] = 16'h3e9b;
mem_array[36527] = 16'heec5;
mem_array[36526] = 16'hbc30;
mem_array[36529] = 16'hbfdb;
mem_array[36528] = 16'h3de2;
mem_array[36531] = 16'h1254;
mem_array[36530] = 16'hbf77;
mem_array[36533] = 16'h3c82;
mem_array[36532] = 16'h3df8;
mem_array[36535] = 16'h8639;
mem_array[36534] = 16'h3df4;
mem_array[36537] = 16'he62f;
mem_array[36536] = 16'hbd01;
mem_array[36539] = 16'hb396;
mem_array[36538] = 16'hbf1a;
mem_array[36541] = 16'ha5f3;
mem_array[36540] = 16'hbd4e;
mem_array[36543] = 16'h4f30;
mem_array[36542] = 16'hbcd7;
mem_array[36545] = 16'he154;
mem_array[36544] = 16'hbde9;
mem_array[36547] = 16'h8a17;
mem_array[36546] = 16'hbee6;
mem_array[36549] = 16'hfbe2;
mem_array[36548] = 16'h3e96;
mem_array[36551] = 16'h49d5;
mem_array[36550] = 16'h3e26;
mem_array[36553] = 16'h9e9c;
mem_array[36552] = 16'hbed8;
mem_array[36555] = 16'h9dac;
mem_array[36554] = 16'h3d85;
mem_array[36557] = 16'h521b;
mem_array[36556] = 16'hbe97;
mem_array[36559] = 16'h78c2;
mem_array[36558] = 16'h3e6a;
mem_array[36561] = 16'h2527;
mem_array[36560] = 16'h3bc4;
mem_array[36563] = 16'h948b;
mem_array[36562] = 16'h3d39;
mem_array[36565] = 16'h1b71;
mem_array[36564] = 16'hbeda;
mem_array[36567] = 16'he779;
mem_array[36566] = 16'h3f2b;
mem_array[36569] = 16'h4b5d;
mem_array[36568] = 16'h3d81;
mem_array[36571] = 16'hf4aa;
mem_array[36570] = 16'hbdb8;
mem_array[36573] = 16'hba88;
mem_array[36572] = 16'hbd35;
mem_array[36575] = 16'ha603;
mem_array[36574] = 16'hbe4d;
mem_array[36577] = 16'hf8d7;
mem_array[36576] = 16'hbef9;
mem_array[36579] = 16'hac53;
mem_array[36578] = 16'h3ea3;
mem_array[36581] = 16'h1fd5;
mem_array[36580] = 16'hbf06;
mem_array[36583] = 16'h0118;
mem_array[36582] = 16'h3e18;
mem_array[36585] = 16'h7845;
mem_array[36584] = 16'hbe00;
mem_array[36587] = 16'h6ec0;
mem_array[36586] = 16'h3e3b;
mem_array[36589] = 16'h1644;
mem_array[36588] = 16'h3cea;
mem_array[36591] = 16'h0533;
mem_array[36590] = 16'hbd35;
mem_array[36593] = 16'h4132;
mem_array[36592] = 16'hbda6;
mem_array[36595] = 16'hcacc;
mem_array[36594] = 16'hbe2b;
mem_array[36597] = 16'hb5c0;
mem_array[36596] = 16'h3e60;
mem_array[36599] = 16'h273d;
mem_array[36598] = 16'hbf82;
mem_array[36601] = 16'hf930;
mem_array[36600] = 16'h3ede;
mem_array[36603] = 16'hde16;
mem_array[36602] = 16'h3e16;
mem_array[36605] = 16'hff68;
mem_array[36604] = 16'h3ec5;
mem_array[36607] = 16'hb26c;
mem_array[36606] = 16'hbe6e;
mem_array[36609] = 16'h95da;
mem_array[36608] = 16'hbde5;
mem_array[36611] = 16'hafbd;
mem_array[36610] = 16'hbf44;
mem_array[36613] = 16'hc302;
mem_array[36612] = 16'hbe9d;
mem_array[36615] = 16'hb315;
mem_array[36614] = 16'hbe99;
mem_array[36617] = 16'h2ce2;
mem_array[36616] = 16'hbf34;
mem_array[36619] = 16'hca47;
mem_array[36618] = 16'hbe18;
mem_array[36621] = 16'h5a11;
mem_array[36620] = 16'hbd8d;
mem_array[36623] = 16'h997b;
mem_array[36622] = 16'hbd0a;
mem_array[36625] = 16'h0b2a;
mem_array[36624] = 16'h3e16;
mem_array[36627] = 16'h1a97;
mem_array[36626] = 16'h3f18;
mem_array[36629] = 16'h0420;
mem_array[36628] = 16'hbe00;
mem_array[36631] = 16'h2a88;
mem_array[36630] = 16'hbe29;
mem_array[36633] = 16'h54ad;
mem_array[36632] = 16'h3f7e;
mem_array[36635] = 16'h0d15;
mem_array[36634] = 16'h3e9c;
mem_array[36637] = 16'h589f;
mem_array[36636] = 16'hbf11;
mem_array[36639] = 16'h6dc2;
mem_array[36638] = 16'hbba6;
mem_array[36641] = 16'hc04c;
mem_array[36640] = 16'h3cf7;
mem_array[36643] = 16'h0d66;
mem_array[36642] = 16'h3d1c;
mem_array[36645] = 16'hd9d2;
mem_array[36644] = 16'hbe13;
mem_array[36647] = 16'haa56;
mem_array[36646] = 16'h3e2c;
mem_array[36649] = 16'h6961;
mem_array[36648] = 16'hbdce;
mem_array[36651] = 16'he431;
mem_array[36650] = 16'hbe88;
mem_array[36653] = 16'hf861;
mem_array[36652] = 16'h3e68;
mem_array[36655] = 16'h85dc;
mem_array[36654] = 16'hbd0c;
mem_array[36657] = 16'h4127;
mem_array[36656] = 16'h3eb3;
mem_array[36659] = 16'hddad;
mem_array[36658] = 16'hbf62;
mem_array[36661] = 16'h544e;
mem_array[36660] = 16'h3ed8;
mem_array[36663] = 16'he4f2;
mem_array[36662] = 16'hbeb9;
mem_array[36665] = 16'h9dff;
mem_array[36664] = 16'h3f4d;
mem_array[36667] = 16'hf904;
mem_array[36666] = 16'hbd10;
mem_array[36669] = 16'h7352;
mem_array[36668] = 16'hbd8d;
mem_array[36671] = 16'h0654;
mem_array[36670] = 16'hbf8c;
mem_array[36673] = 16'hfb5f;
mem_array[36672] = 16'hbe30;
mem_array[36675] = 16'h3b48;
mem_array[36674] = 16'hbebb;
mem_array[36677] = 16'hc46b;
mem_array[36676] = 16'hbf1b;
mem_array[36679] = 16'hc8e6;
mem_array[36678] = 16'h3d1f;
mem_array[36681] = 16'ha30b;
mem_array[36680] = 16'h3ae5;
mem_array[36683] = 16'hb9d5;
mem_array[36682] = 16'h3def;
mem_array[36685] = 16'hca70;
mem_array[36684] = 16'hbefa;
mem_array[36687] = 16'h134f;
mem_array[36686] = 16'h3ec2;
mem_array[36689] = 16'h853c;
mem_array[36688] = 16'hbe63;
mem_array[36691] = 16'hb486;
mem_array[36690] = 16'hbecf;
mem_array[36693] = 16'he45f;
mem_array[36692] = 16'h3ded;
mem_array[36695] = 16'h62ae;
mem_array[36694] = 16'hbe13;
mem_array[36697] = 16'hfb41;
mem_array[36696] = 16'hbf83;
mem_array[36699] = 16'hd493;
mem_array[36698] = 16'h3edf;
mem_array[36701] = 16'h87ee;
mem_array[36700] = 16'h3c10;
mem_array[36703] = 16'h3fc0;
mem_array[36702] = 16'h3ebc;
mem_array[36705] = 16'h8ea1;
mem_array[36704] = 16'h3eeb;
mem_array[36707] = 16'h0f7f;
mem_array[36706] = 16'hbec2;
mem_array[36709] = 16'ha089;
mem_array[36708] = 16'hbe80;
mem_array[36711] = 16'h2f60;
mem_array[36710] = 16'hbf35;
mem_array[36713] = 16'h507b;
mem_array[36712] = 16'h3f21;
mem_array[36715] = 16'h41f2;
mem_array[36714] = 16'h3f0b;
mem_array[36717] = 16'hccc5;
mem_array[36716] = 16'hbdbd;
mem_array[36719] = 16'hfbfd;
mem_array[36718] = 16'hbe90;
mem_array[36721] = 16'h78cf;
mem_array[36720] = 16'h3ee6;
mem_array[36723] = 16'hd359;
mem_array[36722] = 16'h3f28;
mem_array[36725] = 16'h4b84;
mem_array[36724] = 16'h3ebd;
mem_array[36727] = 16'h9317;
mem_array[36726] = 16'hbdaf;
mem_array[36729] = 16'h03ba;
mem_array[36728] = 16'h3ec0;
mem_array[36731] = 16'h9ea0;
mem_array[36730] = 16'hbe23;
mem_array[36733] = 16'ha6e1;
mem_array[36732] = 16'hbf10;
mem_array[36735] = 16'hb107;
mem_array[36734] = 16'hbef9;
mem_array[36737] = 16'h808f;
mem_array[36736] = 16'hbebf;
mem_array[36739] = 16'h8414;
mem_array[36738] = 16'h3e2f;
mem_array[36741] = 16'h366d;
mem_array[36740] = 16'h3c4c;
mem_array[36743] = 16'h3265;
mem_array[36742] = 16'h3d76;
mem_array[36745] = 16'h9785;
mem_array[36744] = 16'hbf42;
mem_array[36747] = 16'hfd50;
mem_array[36746] = 16'h3f1a;
mem_array[36749] = 16'h479f;
mem_array[36748] = 16'h3f1c;
mem_array[36751] = 16'h77db;
mem_array[36750] = 16'hbe80;
mem_array[36753] = 16'hcfcd;
mem_array[36752] = 16'h3f1e;
mem_array[36755] = 16'hf171;
mem_array[36754] = 16'h3e99;
mem_array[36757] = 16'h9be1;
mem_array[36756] = 16'h3f05;
mem_array[36759] = 16'h844b;
mem_array[36758] = 16'h3f49;
mem_array[36761] = 16'hc9ac;
mem_array[36760] = 16'hbefd;
mem_array[36763] = 16'he9e5;
mem_array[36762] = 16'hbb8f;
mem_array[36765] = 16'hd0a8;
mem_array[36764] = 16'hbfaa;
mem_array[36767] = 16'h61a0;
mem_array[36766] = 16'hbee9;
mem_array[36769] = 16'h91a6;
mem_array[36768] = 16'h3ef6;
mem_array[36771] = 16'h774f;
mem_array[36770] = 16'hbd8a;
mem_array[36773] = 16'h754c;
mem_array[36772] = 16'h3e97;
mem_array[36775] = 16'h6b10;
mem_array[36774] = 16'hbe3f;
mem_array[36777] = 16'h29fe;
mem_array[36776] = 16'h3e97;
mem_array[36779] = 16'hc807;
mem_array[36778] = 16'hbf65;
mem_array[36781] = 16'h65a0;
mem_array[36780] = 16'h3f35;
mem_array[36783] = 16'h3007;
mem_array[36782] = 16'hbe20;
mem_array[36785] = 16'hb347;
mem_array[36784] = 16'h402f;
mem_array[36787] = 16'hd9d3;
mem_array[36786] = 16'hbe49;
mem_array[36789] = 16'hbca6;
mem_array[36788] = 16'hbdba;
mem_array[36791] = 16'h04f4;
mem_array[36790] = 16'hbe27;
mem_array[36793] = 16'h6f15;
mem_array[36792] = 16'h3f15;
mem_array[36795] = 16'h880d;
mem_array[36794] = 16'hbe8d;
mem_array[36797] = 16'h9f9c;
mem_array[36796] = 16'h3e83;
mem_array[36799] = 16'h99a3;
mem_array[36798] = 16'h3f7e;
mem_array[36801] = 16'h3ded;
mem_array[36800] = 16'hbd00;
mem_array[36803] = 16'hb496;
mem_array[36802] = 16'h3d76;
mem_array[36805] = 16'h3511;
mem_array[36804] = 16'h3d27;
mem_array[36807] = 16'h7030;
mem_array[36806] = 16'h3f14;
mem_array[36809] = 16'h5fe4;
mem_array[36808] = 16'h3f69;
mem_array[36811] = 16'hffa6;
mem_array[36810] = 16'hbf8a;
mem_array[36813] = 16'h33a5;
mem_array[36812] = 16'h3fdb;
mem_array[36815] = 16'hb88e;
mem_array[36814] = 16'hbe8d;
mem_array[36817] = 16'h4868;
mem_array[36816] = 16'h3f4c;
mem_array[36819] = 16'h0db8;
mem_array[36818] = 16'h3e4b;
mem_array[36821] = 16'he12c;
mem_array[36820] = 16'hbe8b;
mem_array[36823] = 16'h2a17;
mem_array[36822] = 16'h3d62;
mem_array[36825] = 16'h42e2;
mem_array[36824] = 16'hbec3;
mem_array[36827] = 16'hee48;
mem_array[36826] = 16'h3e3b;
mem_array[36829] = 16'he725;
mem_array[36828] = 16'h3f69;
mem_array[36831] = 16'h84bb;
mem_array[36830] = 16'h3d38;
mem_array[36833] = 16'hc08f;
mem_array[36832] = 16'h3ed9;
mem_array[36835] = 16'h1f8f;
mem_array[36834] = 16'hbf38;
mem_array[36837] = 16'h88e0;
mem_array[36836] = 16'h3ed5;
mem_array[36839] = 16'h7d0b;
mem_array[36838] = 16'hbf2a;
mem_array[36841] = 16'h2493;
mem_array[36840] = 16'h3f66;
mem_array[36843] = 16'h1bed;
mem_array[36842] = 16'h3d83;
mem_array[36845] = 16'h87e3;
mem_array[36844] = 16'h3f93;
mem_array[36847] = 16'h7a68;
mem_array[36846] = 16'h3fcd;
mem_array[36849] = 16'h0bc2;
mem_array[36848] = 16'h3b69;
mem_array[36851] = 16'h0d1d;
mem_array[36850] = 16'h3eee;
mem_array[36853] = 16'h3233;
mem_array[36852] = 16'hbc87;
mem_array[36855] = 16'haf26;
mem_array[36854] = 16'hbee8;
mem_array[36857] = 16'h2248;
mem_array[36856] = 16'h3eab;
mem_array[36859] = 16'h6be0;
mem_array[36858] = 16'h3f34;
mem_array[36861] = 16'h73b7;
mem_array[36860] = 16'h3d2a;
mem_array[36863] = 16'h660d;
mem_array[36862] = 16'hb9de;
mem_array[36865] = 16'h6cab;
mem_array[36864] = 16'h3f43;
mem_array[36867] = 16'hf227;
mem_array[36866] = 16'hbeef;
mem_array[36869] = 16'h019a;
mem_array[36868] = 16'h3e2a;
mem_array[36871] = 16'h0e8f;
mem_array[36870] = 16'hbf3b;
mem_array[36873] = 16'h9b02;
mem_array[36872] = 16'h3f92;
mem_array[36875] = 16'hf4fc;
mem_array[36874] = 16'h3d20;
mem_array[36877] = 16'h0753;
mem_array[36876] = 16'hbf92;
mem_array[36879] = 16'he3b5;
mem_array[36878] = 16'hbed5;
mem_array[36881] = 16'h262f;
mem_array[36880] = 16'h3b8c;
mem_array[36883] = 16'h6982;
mem_array[36882] = 16'h3f38;
mem_array[36885] = 16'h2270;
mem_array[36884] = 16'hbdbe;
mem_array[36887] = 16'hcaf2;
mem_array[36886] = 16'h3efc;
mem_array[36889] = 16'h59f2;
mem_array[36888] = 16'h3ec0;
mem_array[36891] = 16'h9df2;
mem_array[36890] = 16'h3d88;
mem_array[36893] = 16'ha3b0;
mem_array[36892] = 16'h3e13;
mem_array[36895] = 16'h62d3;
mem_array[36894] = 16'hbeba;
mem_array[36897] = 16'h5134;
mem_array[36896] = 16'hbe05;
mem_array[36899] = 16'h2f97;
mem_array[36898] = 16'h3ee6;
mem_array[36901] = 16'h0b6c;
mem_array[36900] = 16'h3de6;
mem_array[36903] = 16'h712d;
mem_array[36902] = 16'hbdbc;
mem_array[36905] = 16'hb8ed;
mem_array[36904] = 16'hbd49;
mem_array[36907] = 16'h0ba8;
mem_array[36906] = 16'hbd66;
mem_array[36909] = 16'h0ba6;
mem_array[36908] = 16'h3db3;
mem_array[36911] = 16'h55be;
mem_array[36910] = 16'hbd44;
mem_array[36913] = 16'hf3bb;
mem_array[36912] = 16'hbd96;
mem_array[36915] = 16'h2d93;
mem_array[36914] = 16'hbd5b;
mem_array[36917] = 16'hab56;
mem_array[36916] = 16'h3d0d;
mem_array[36919] = 16'h6041;
mem_array[36918] = 16'h3d2f;
mem_array[36921] = 16'h8d3e;
mem_array[36920] = 16'h3ce6;
mem_array[36923] = 16'h1340;
mem_array[36922] = 16'hbd4f;
mem_array[36925] = 16'heefc;
mem_array[36924] = 16'h3cdb;
mem_array[36927] = 16'hff66;
mem_array[36926] = 16'h3c1c;
mem_array[36929] = 16'h4df1;
mem_array[36928] = 16'hbd3e;
mem_array[36931] = 16'h5c04;
mem_array[36930] = 16'h3d09;
mem_array[36933] = 16'ha282;
mem_array[36932] = 16'h3bad;
mem_array[36935] = 16'h2ddf;
mem_array[36934] = 16'hbbb9;
mem_array[36937] = 16'h1432;
mem_array[36936] = 16'h3cb2;
mem_array[36939] = 16'h4721;
mem_array[36938] = 16'h3d0c;
mem_array[36941] = 16'h6779;
mem_array[36940] = 16'hbda3;
mem_array[36943] = 16'h6dcc;
mem_array[36942] = 16'h3c6c;
mem_array[36945] = 16'h11f3;
mem_array[36944] = 16'hbc94;
mem_array[36947] = 16'h5c42;
mem_array[36946] = 16'h3c08;
mem_array[36949] = 16'he981;
mem_array[36948] = 16'hbce5;
mem_array[36951] = 16'h1a66;
mem_array[36950] = 16'h3d64;
mem_array[36953] = 16'h97ba;
mem_array[36952] = 16'hbd9c;
mem_array[36955] = 16'h0ad4;
mem_array[36954] = 16'h3d91;
mem_array[36957] = 16'h302b;
mem_array[36956] = 16'h3d1b;
mem_array[36959] = 16'h3a5a;
mem_array[36958] = 16'h3ad9;
mem_array[36961] = 16'hccdf;
mem_array[36960] = 16'hbcf5;
mem_array[36963] = 16'hc007;
mem_array[36962] = 16'h3d90;
mem_array[36965] = 16'h7d84;
mem_array[36964] = 16'h3d32;
mem_array[36967] = 16'hdd9c;
mem_array[36966] = 16'hbd9e;
mem_array[36969] = 16'h563a;
mem_array[36968] = 16'h3d9e;
mem_array[36971] = 16'h34b9;
mem_array[36970] = 16'hbd63;
mem_array[36973] = 16'hf37b;
mem_array[36972] = 16'h3d94;
mem_array[36975] = 16'h2284;
mem_array[36974] = 16'h3d0a;
mem_array[36977] = 16'h71be;
mem_array[36976] = 16'h3d81;
mem_array[36979] = 16'ha9c8;
mem_array[36978] = 16'h3dd3;
mem_array[36981] = 16'haa96;
mem_array[36980] = 16'h3dbe;
mem_array[36983] = 16'h61e6;
mem_array[36982] = 16'h3c85;
mem_array[36985] = 16'hec6d;
mem_array[36984] = 16'h3dcc;
mem_array[36987] = 16'h2bfd;
mem_array[36986] = 16'hbbba;
mem_array[36989] = 16'h9fb7;
mem_array[36988] = 16'h3be3;
mem_array[36991] = 16'h4d4b;
mem_array[36990] = 16'h3dd1;
mem_array[36993] = 16'h8b6e;
mem_array[36992] = 16'hbd91;
mem_array[36995] = 16'h9d68;
mem_array[36994] = 16'h3b5f;
mem_array[36997] = 16'hcefd;
mem_array[36996] = 16'h3c46;
mem_array[36999] = 16'hcfeb;
mem_array[36998] = 16'hbc93;
mem_array[37001] = 16'he8a2;
mem_array[37000] = 16'h3db9;
mem_array[37003] = 16'h3456;
mem_array[37002] = 16'h3db2;
mem_array[37005] = 16'h82c9;
mem_array[37004] = 16'hbdab;
mem_array[37007] = 16'heb9f;
mem_array[37006] = 16'hbca3;
mem_array[37009] = 16'hc946;
mem_array[37008] = 16'hbcc6;
mem_array[37011] = 16'ha75b;
mem_array[37010] = 16'hbc15;
mem_array[37013] = 16'hdd7b;
mem_array[37012] = 16'h3c1f;
mem_array[37015] = 16'hbb6f;
mem_array[37014] = 16'h3c8d;
mem_array[37017] = 16'h854f;
mem_array[37016] = 16'hbd88;
mem_array[37019] = 16'hf6a3;
mem_array[37018] = 16'h3d32;
mem_array[37021] = 16'h23c2;
mem_array[37020] = 16'hbd81;
mem_array[37023] = 16'h91c2;
mem_array[37022] = 16'h3dc9;
mem_array[37025] = 16'h3b20;
mem_array[37024] = 16'h3da1;
mem_array[37027] = 16'h5381;
mem_array[37026] = 16'hbd34;
mem_array[37029] = 16'h3269;
mem_array[37028] = 16'h3b98;
mem_array[37031] = 16'hb025;
mem_array[37030] = 16'hbded;
mem_array[37033] = 16'hb62a;
mem_array[37032] = 16'h3e83;
mem_array[37035] = 16'hc5ac;
mem_array[37034] = 16'h3c56;
mem_array[37037] = 16'he1b4;
mem_array[37036] = 16'h3cc2;
mem_array[37039] = 16'h6e07;
mem_array[37038] = 16'h3cce;
mem_array[37041] = 16'h3938;
mem_array[37040] = 16'hbd9e;
mem_array[37043] = 16'h359f;
mem_array[37042] = 16'hbd9d;
mem_array[37045] = 16'had8c;
mem_array[37044] = 16'hbc01;
mem_array[37047] = 16'h1425;
mem_array[37046] = 16'hbddf;
mem_array[37049] = 16'h0a8d;
mem_array[37048] = 16'h3dc6;
mem_array[37051] = 16'h55c3;
mem_array[37050] = 16'h3e5a;
mem_array[37053] = 16'hb853;
mem_array[37052] = 16'h3d52;
mem_array[37055] = 16'h50bc;
mem_array[37054] = 16'h3d87;
mem_array[37057] = 16'h78a9;
mem_array[37056] = 16'h3ccf;
mem_array[37059] = 16'hc536;
mem_array[37058] = 16'hbc00;
mem_array[37061] = 16'hb772;
mem_array[37060] = 16'h3d4f;
mem_array[37063] = 16'h90fe;
mem_array[37062] = 16'h3edc;
mem_array[37065] = 16'h969b;
mem_array[37064] = 16'h3cb1;
mem_array[37067] = 16'hde4b;
mem_array[37066] = 16'hbd9f;
mem_array[37069] = 16'he086;
mem_array[37068] = 16'h3e82;
mem_array[37071] = 16'hccb7;
mem_array[37070] = 16'h3d5d;
mem_array[37073] = 16'h2f0b;
mem_array[37072] = 16'h3e12;
mem_array[37075] = 16'hc055;
mem_array[37074] = 16'hbd8d;
mem_array[37077] = 16'h5fa6;
mem_array[37076] = 16'h3c61;
mem_array[37079] = 16'h0067;
mem_array[37078] = 16'h3d71;
mem_array[37081] = 16'h97a7;
mem_array[37080] = 16'h3e00;
mem_array[37083] = 16'h2390;
mem_array[37082] = 16'h3e40;
mem_array[37085] = 16'hecb9;
mem_array[37084] = 16'h3fc0;
mem_array[37087] = 16'h916e;
mem_array[37086] = 16'h3d5c;
mem_array[37089] = 16'h8e66;
mem_array[37088] = 16'hbdfa;
mem_array[37091] = 16'h8816;
mem_array[37090] = 16'hbd97;
mem_array[37093] = 16'hbe2c;
mem_array[37092] = 16'hbd87;
mem_array[37095] = 16'hb3c3;
mem_array[37094] = 16'hbe6c;
mem_array[37097] = 16'ha04c;
mem_array[37096] = 16'h3eb4;
mem_array[37099] = 16'hb0eb;
mem_array[37098] = 16'h3aff;
mem_array[37101] = 16'h7b09;
mem_array[37100] = 16'h3b82;
mem_array[37103] = 16'he6dd;
mem_array[37102] = 16'h3cd5;
mem_array[37105] = 16'h2346;
mem_array[37104] = 16'hbec1;
mem_array[37107] = 16'h33da;
mem_array[37106] = 16'h3f2c;
mem_array[37109] = 16'hc0cf;
mem_array[37108] = 16'h3ed9;
mem_array[37111] = 16'h56cd;
mem_array[37110] = 16'hbe10;
mem_array[37113] = 16'h7a47;
mem_array[37112] = 16'hbe3b;
mem_array[37115] = 16'ha9e7;
mem_array[37114] = 16'h3e0d;
mem_array[37117] = 16'h9704;
mem_array[37116] = 16'hbe4b;
mem_array[37119] = 16'h5e16;
mem_array[37118] = 16'hbe8c;
mem_array[37121] = 16'h5705;
mem_array[37120] = 16'hbdbc;
mem_array[37123] = 16'h0e83;
mem_array[37122] = 16'h3ee7;
mem_array[37125] = 16'hb11f;
mem_array[37124] = 16'hbc7c;
mem_array[37127] = 16'h65b4;
mem_array[37126] = 16'hbd6b;
mem_array[37129] = 16'hf6cc;
mem_array[37128] = 16'hbb61;
mem_array[37131] = 16'h2bdb;
mem_array[37130] = 16'hbd33;
mem_array[37133] = 16'h9bfe;
mem_array[37132] = 16'hbe81;
mem_array[37135] = 16'h5c7e;
mem_array[37134] = 16'h3f0a;
mem_array[37137] = 16'h8a8e;
mem_array[37136] = 16'hbeb9;
mem_array[37139] = 16'h1e2e;
mem_array[37138] = 16'hbe00;
mem_array[37141] = 16'h8563;
mem_array[37140] = 16'hbdf4;
mem_array[37143] = 16'hcec7;
mem_array[37142] = 16'hbf5e;
mem_array[37145] = 16'h19a2;
mem_array[37144] = 16'h3ea7;
mem_array[37147] = 16'h1120;
mem_array[37146] = 16'h3de3;
mem_array[37149] = 16'h50d6;
mem_array[37148] = 16'h3eda;
mem_array[37151] = 16'h19b7;
mem_array[37150] = 16'h3e0a;
mem_array[37153] = 16'hfd2f;
mem_array[37152] = 16'hbe00;
mem_array[37155] = 16'h5225;
mem_array[37154] = 16'hbdad;
mem_array[37157] = 16'ha7fd;
mem_array[37156] = 16'h3e6e;
mem_array[37159] = 16'h7581;
mem_array[37158] = 16'hbda8;
mem_array[37161] = 16'h8ca2;
mem_array[37160] = 16'hbdbc;
mem_array[37163] = 16'h4ea8;
mem_array[37162] = 16'hbdb4;
mem_array[37165] = 16'hbce5;
mem_array[37164] = 16'h3e6b;
mem_array[37167] = 16'h038b;
mem_array[37166] = 16'h3f8a;
mem_array[37169] = 16'h3ba3;
mem_array[37168] = 16'h3d0e;
mem_array[37171] = 16'he42d;
mem_array[37170] = 16'hbeeb;
mem_array[37173] = 16'h5409;
mem_array[37172] = 16'h3fa5;
mem_array[37175] = 16'h41dd;
mem_array[37174] = 16'hbea9;
mem_array[37177] = 16'h2d47;
mem_array[37176] = 16'hbec2;
mem_array[37179] = 16'h1c42;
mem_array[37178] = 16'hbfc5;
mem_array[37181] = 16'h8f7c;
mem_array[37180] = 16'hbee9;
mem_array[37183] = 16'hbc2b;
mem_array[37182] = 16'h3df7;
mem_array[37185] = 16'h04ff;
mem_array[37184] = 16'hbbcb;
mem_array[37187] = 16'h6afa;
mem_array[37186] = 16'h3bad;
mem_array[37189] = 16'hab67;
mem_array[37188] = 16'h3e04;
mem_array[37191] = 16'h88de;
mem_array[37190] = 16'hbf0b;
mem_array[37193] = 16'h8730;
mem_array[37192] = 16'h3de7;
mem_array[37195] = 16'h5d95;
mem_array[37194] = 16'hbee5;
mem_array[37197] = 16'h765c;
mem_array[37196] = 16'h3cee;
mem_array[37199] = 16'h1a4c;
mem_array[37198] = 16'hbe6a;
mem_array[37201] = 16'h6521;
mem_array[37200] = 16'h3f54;
mem_array[37203] = 16'h99aa;
mem_array[37202] = 16'hbf4e;
mem_array[37205] = 16'h0cad;
mem_array[37204] = 16'h3dc6;
mem_array[37207] = 16'h3af7;
mem_array[37206] = 16'hbec1;
mem_array[37209] = 16'h8ef6;
mem_array[37208] = 16'h3f1c;
mem_array[37211] = 16'h3a16;
mem_array[37210] = 16'hbee1;
mem_array[37213] = 16'h4319;
mem_array[37212] = 16'h3e4d;
mem_array[37215] = 16'hbd31;
mem_array[37214] = 16'hbdeb;
mem_array[37217] = 16'hd011;
mem_array[37216] = 16'h3e97;
mem_array[37219] = 16'h9850;
mem_array[37218] = 16'hbe1e;
mem_array[37221] = 16'h9a21;
mem_array[37220] = 16'hbbcf;
mem_array[37223] = 16'h4509;
mem_array[37222] = 16'hbd83;
mem_array[37225] = 16'hd27b;
mem_array[37224] = 16'hbe9e;
mem_array[37227] = 16'h147b;
mem_array[37226] = 16'hbe6f;
mem_array[37229] = 16'h0099;
mem_array[37228] = 16'h3bda;
mem_array[37231] = 16'h2da9;
mem_array[37230] = 16'h3d5c;
mem_array[37233] = 16'hf8e5;
mem_array[37232] = 16'h3db8;
mem_array[37235] = 16'h004b;
mem_array[37234] = 16'h3f4b;
mem_array[37237] = 16'he6b8;
mem_array[37236] = 16'hbfa8;
mem_array[37239] = 16'hfd83;
mem_array[37238] = 16'hbfd3;
mem_array[37241] = 16'h9136;
mem_array[37240] = 16'h3e3b;
mem_array[37243] = 16'hb1f5;
mem_array[37242] = 16'hbda3;
mem_array[37245] = 16'hc377;
mem_array[37244] = 16'hbe06;
mem_array[37247] = 16'h7292;
mem_array[37246] = 16'h3ecc;
mem_array[37249] = 16'hc266;
mem_array[37248] = 16'hbe31;
mem_array[37251] = 16'h0065;
mem_array[37250] = 16'hbeb1;
mem_array[37253] = 16'hafcd;
mem_array[37252] = 16'h3cc2;
mem_array[37255] = 16'h768f;
mem_array[37254] = 16'h3e87;
mem_array[37257] = 16'ha5d7;
mem_array[37256] = 16'hbeb5;
mem_array[37259] = 16'h0a45;
mem_array[37258] = 16'hbfd0;
mem_array[37261] = 16'h1070;
mem_array[37260] = 16'h3eee;
mem_array[37263] = 16'he444;
mem_array[37262] = 16'hbe19;
mem_array[37265] = 16'h57f9;
mem_array[37264] = 16'hbf22;
mem_array[37267] = 16'he541;
mem_array[37266] = 16'h3f38;
mem_array[37269] = 16'he340;
mem_array[37268] = 16'hbe1f;
mem_array[37271] = 16'hbbfd;
mem_array[37270] = 16'h3ed3;
mem_array[37273] = 16'h2264;
mem_array[37272] = 16'h3d13;
mem_array[37275] = 16'h6021;
mem_array[37274] = 16'hbeb5;
mem_array[37277] = 16'h3a7e;
mem_array[37276] = 16'h3d5d;
mem_array[37279] = 16'hdec0;
mem_array[37278] = 16'hbee8;
mem_array[37281] = 16'h5a7d;
mem_array[37280] = 16'hbd02;
mem_array[37283] = 16'he588;
mem_array[37282] = 16'hbd95;
mem_array[37285] = 16'hc644;
mem_array[37284] = 16'h3d6b;
mem_array[37287] = 16'h7c09;
mem_array[37286] = 16'hbe83;
mem_array[37289] = 16'h0c52;
mem_array[37288] = 16'h3e90;
mem_array[37291] = 16'h4ad2;
mem_array[37290] = 16'h3e60;
mem_array[37293] = 16'haa91;
mem_array[37292] = 16'hbe05;
mem_array[37295] = 16'h3d00;
mem_array[37294] = 16'h3ed0;
mem_array[37297] = 16'hc513;
mem_array[37296] = 16'hbfa4;
mem_array[37299] = 16'h997d;
mem_array[37298] = 16'hbe58;
mem_array[37301] = 16'h0e08;
mem_array[37300] = 16'hbf54;
mem_array[37303] = 16'h531c;
mem_array[37302] = 16'hbca1;
mem_array[37305] = 16'h4910;
mem_array[37304] = 16'hbf2e;
mem_array[37307] = 16'h62ed;
mem_array[37306] = 16'hbea0;
mem_array[37309] = 16'hdff9;
mem_array[37308] = 16'h3e64;
mem_array[37311] = 16'hf23e;
mem_array[37310] = 16'h3d69;
mem_array[37313] = 16'h8f91;
mem_array[37312] = 16'hbd01;
mem_array[37315] = 16'hccb5;
mem_array[37314] = 16'h3e5c;
mem_array[37317] = 16'h402f;
mem_array[37316] = 16'h3e4e;
mem_array[37319] = 16'h33c9;
mem_array[37318] = 16'hbfbc;
mem_array[37321] = 16'hcbe2;
mem_array[37320] = 16'h3dae;
mem_array[37323] = 16'h27e2;
mem_array[37322] = 16'hbf72;
mem_array[37325] = 16'hf37a;
mem_array[37324] = 16'hbe96;
mem_array[37327] = 16'h8ed3;
mem_array[37326] = 16'h3db1;
mem_array[37329] = 16'h2d9e;
mem_array[37328] = 16'hbd77;
mem_array[37331] = 16'h3b26;
mem_array[37330] = 16'hbe76;
mem_array[37333] = 16'hf5bc;
mem_array[37332] = 16'h3ec5;
mem_array[37335] = 16'h9f7b;
mem_array[37334] = 16'hbefe;
mem_array[37337] = 16'hfd61;
mem_array[37336] = 16'h3def;
mem_array[37339] = 16'hdb8b;
mem_array[37338] = 16'h3d04;
mem_array[37341] = 16'h20bf;
mem_array[37340] = 16'hbb8f;
mem_array[37343] = 16'h1c65;
mem_array[37342] = 16'h3c84;
mem_array[37345] = 16'h22f9;
mem_array[37344] = 16'h3f16;
mem_array[37347] = 16'hbc71;
mem_array[37346] = 16'hbe39;
mem_array[37349] = 16'hcff1;
mem_array[37348] = 16'h3e46;
mem_array[37351] = 16'h23a0;
mem_array[37350] = 16'h3eb1;
mem_array[37353] = 16'h9c8e;
mem_array[37352] = 16'h3e4a;
mem_array[37355] = 16'hc047;
mem_array[37354] = 16'h3dac;
mem_array[37357] = 16'hefc2;
mem_array[37356] = 16'hbf81;
mem_array[37359] = 16'hc5fc;
mem_array[37358] = 16'hbf5e;
mem_array[37361] = 16'h1f86;
mem_array[37360] = 16'hbe69;
mem_array[37363] = 16'h87ec;
mem_array[37362] = 16'h3ca7;
mem_array[37365] = 16'hdc89;
mem_array[37364] = 16'hbfe0;
mem_array[37367] = 16'h1437;
mem_array[37366] = 16'h3de7;
mem_array[37369] = 16'h5f12;
mem_array[37368] = 16'hbebb;
mem_array[37371] = 16'h3900;
mem_array[37370] = 16'hbced;
mem_array[37373] = 16'h6818;
mem_array[37372] = 16'hbe04;
mem_array[37375] = 16'h84af;
mem_array[37374] = 16'h3c9b;
mem_array[37377] = 16'hfb09;
mem_array[37376] = 16'h3ea1;
mem_array[37379] = 16'h99d0;
mem_array[37378] = 16'hbf8d;
mem_array[37381] = 16'h8785;
mem_array[37380] = 16'hbe12;
mem_array[37383] = 16'h285d;
mem_array[37382] = 16'hbe0e;
mem_array[37385] = 16'hf434;
mem_array[37384] = 16'h3e07;
mem_array[37387] = 16'h75f3;
mem_array[37386] = 16'h3e3d;
mem_array[37389] = 16'heefd;
mem_array[37388] = 16'h3e5f;
mem_array[37391] = 16'h60ca;
mem_array[37390] = 16'h3d15;
mem_array[37393] = 16'hf68e;
mem_array[37392] = 16'h3eab;
mem_array[37395] = 16'h1448;
mem_array[37394] = 16'hbe0e;
mem_array[37397] = 16'h27a1;
mem_array[37396] = 16'hbdc2;
mem_array[37399] = 16'hc0aa;
mem_array[37398] = 16'h3e75;
mem_array[37401] = 16'h843d;
mem_array[37400] = 16'hbd1f;
mem_array[37403] = 16'h3c18;
mem_array[37402] = 16'hbc91;
mem_array[37405] = 16'ha448;
mem_array[37404] = 16'h3e86;
mem_array[37407] = 16'he1fc;
mem_array[37406] = 16'hbe79;
mem_array[37409] = 16'h9be5;
mem_array[37408] = 16'h3d16;
mem_array[37411] = 16'h227a;
mem_array[37410] = 16'h3e5e;
mem_array[37413] = 16'h1ed6;
mem_array[37412] = 16'h3e1d;
mem_array[37415] = 16'h0aab;
mem_array[37414] = 16'hbe0f;
mem_array[37417] = 16'ha3ea;
mem_array[37416] = 16'hbfa1;
mem_array[37419] = 16'h05ea;
mem_array[37418] = 16'hbfa9;
mem_array[37421] = 16'h7bf2;
mem_array[37420] = 16'hbefe;
mem_array[37423] = 16'h63f2;
mem_array[37422] = 16'hbe30;
mem_array[37425] = 16'h09c6;
mem_array[37424] = 16'hbe35;
mem_array[37427] = 16'h88e6;
mem_array[37426] = 16'h3e09;
mem_array[37429] = 16'h7c96;
mem_array[37428] = 16'hbafd;
mem_array[37431] = 16'h32b6;
mem_array[37430] = 16'h3de9;
mem_array[37433] = 16'h9563;
mem_array[37432] = 16'hbe5c;
mem_array[37435] = 16'h3fc0;
mem_array[37434] = 16'hbef0;
mem_array[37437] = 16'hcb90;
mem_array[37436] = 16'h3d92;
mem_array[37439] = 16'h55f3;
mem_array[37438] = 16'hbf99;
mem_array[37441] = 16'ha86d;
mem_array[37440] = 16'h3e15;
mem_array[37443] = 16'h65f0;
mem_array[37442] = 16'h3ee6;
mem_array[37445] = 16'h7710;
mem_array[37444] = 16'h3e25;
mem_array[37447] = 16'h882f;
mem_array[37446] = 16'h3e3f;
mem_array[37449] = 16'hd83c;
mem_array[37448] = 16'h3e17;
mem_array[37451] = 16'h27ba;
mem_array[37450] = 16'hbd80;
mem_array[37453] = 16'hb0a1;
mem_array[37452] = 16'hbe4d;
mem_array[37455] = 16'h1922;
mem_array[37454] = 16'hbe76;
mem_array[37457] = 16'hb9ac;
mem_array[37456] = 16'hbd30;
mem_array[37459] = 16'h95f8;
mem_array[37458] = 16'h3e2d;
mem_array[37461] = 16'h000c;
mem_array[37460] = 16'h3aeb;
mem_array[37463] = 16'hc08e;
mem_array[37462] = 16'hbd23;
mem_array[37465] = 16'h5d04;
mem_array[37464] = 16'h3cfa;
mem_array[37467] = 16'h6027;
mem_array[37466] = 16'hbe53;
mem_array[37469] = 16'hb1a7;
mem_array[37468] = 16'h3eab;
mem_array[37471] = 16'h5f6b;
mem_array[37470] = 16'h3ce4;
mem_array[37473] = 16'h02e9;
mem_array[37472] = 16'h3d52;
mem_array[37475] = 16'h47e9;
mem_array[37474] = 16'hbe68;
mem_array[37477] = 16'h8649;
mem_array[37476] = 16'hbe02;
mem_array[37479] = 16'h85cc;
mem_array[37478] = 16'hbfd8;
mem_array[37481] = 16'h1279;
mem_array[37480] = 16'hbe2f;
mem_array[37483] = 16'h3608;
mem_array[37482] = 16'h3e11;
mem_array[37485] = 16'h6571;
mem_array[37484] = 16'hbe9d;
mem_array[37487] = 16'h45ad;
mem_array[37486] = 16'hbe5c;
mem_array[37489] = 16'h8db5;
mem_array[37488] = 16'h3d65;
mem_array[37491] = 16'h56eb;
mem_array[37490] = 16'h3e31;
mem_array[37493] = 16'h26a8;
mem_array[37492] = 16'hbd89;
mem_array[37495] = 16'hc55c;
mem_array[37494] = 16'hbd96;
mem_array[37497] = 16'h235d;
mem_array[37496] = 16'h3e54;
mem_array[37499] = 16'h41fc;
mem_array[37498] = 16'hbe99;
mem_array[37501] = 16'hcc8f;
mem_array[37500] = 16'hbd46;
mem_array[37503] = 16'h565a;
mem_array[37502] = 16'h3e90;
mem_array[37505] = 16'h1d66;
mem_array[37504] = 16'hbd2b;
mem_array[37507] = 16'heb23;
mem_array[37506] = 16'h3cee;
mem_array[37509] = 16'he238;
mem_array[37508] = 16'h3e1e;
mem_array[37511] = 16'h7653;
mem_array[37510] = 16'hbdd8;
mem_array[37513] = 16'h4e73;
mem_array[37512] = 16'h3d67;
mem_array[37515] = 16'h523e;
mem_array[37514] = 16'hbe02;
mem_array[37517] = 16'h24f6;
mem_array[37516] = 16'h3ce1;
mem_array[37519] = 16'h72c6;
mem_array[37518] = 16'hbdb6;
mem_array[37521] = 16'hea15;
mem_array[37520] = 16'hbd67;
mem_array[37523] = 16'hac33;
mem_array[37522] = 16'h3da1;
mem_array[37525] = 16'h9aad;
mem_array[37524] = 16'h3e00;
mem_array[37527] = 16'h438d;
mem_array[37526] = 16'h3d48;
mem_array[37529] = 16'hf2c3;
mem_array[37528] = 16'h3e6a;
mem_array[37531] = 16'hbc8c;
mem_array[37530] = 16'h3d81;
mem_array[37533] = 16'h5d3a;
mem_array[37532] = 16'hbdb5;
mem_array[37535] = 16'h0482;
mem_array[37534] = 16'hbd9d;
mem_array[37537] = 16'h445b;
mem_array[37536] = 16'h3ce8;
mem_array[37539] = 16'h6688;
mem_array[37538] = 16'hbfcd;
mem_array[37541] = 16'h7771;
mem_array[37540] = 16'hbe46;
mem_array[37543] = 16'h2721;
mem_array[37542] = 16'h3eb8;
mem_array[37545] = 16'h796c;
mem_array[37544] = 16'h3d9c;
mem_array[37547] = 16'hf953;
mem_array[37546] = 16'hbe8f;
mem_array[37549] = 16'h4dda;
mem_array[37548] = 16'hbe28;
mem_array[37551] = 16'h0301;
mem_array[37550] = 16'h3e96;
mem_array[37553] = 16'h4ae5;
mem_array[37552] = 16'h3e38;
mem_array[37555] = 16'h0c3e;
mem_array[37554] = 16'h3daa;
mem_array[37557] = 16'had11;
mem_array[37556] = 16'hbdc2;
mem_array[37559] = 16'h3a6b;
mem_array[37558] = 16'h3d45;
mem_array[37561] = 16'h70b4;
mem_array[37560] = 16'hbe36;
mem_array[37563] = 16'h1709;
mem_array[37562] = 16'hbe82;
mem_array[37565] = 16'hde9c;
mem_array[37564] = 16'h3d85;
mem_array[37567] = 16'hc1b4;
mem_array[37566] = 16'h3e4f;
mem_array[37569] = 16'he625;
mem_array[37568] = 16'h3d6b;
mem_array[37571] = 16'h58f4;
mem_array[37570] = 16'hbebd;
mem_array[37573] = 16'h27bf;
mem_array[37572] = 16'h3df4;
mem_array[37575] = 16'hdf86;
mem_array[37574] = 16'h3cac;
mem_array[37577] = 16'hf0fa;
mem_array[37576] = 16'hbefa;
mem_array[37579] = 16'h58b4;
mem_array[37578] = 16'h3e4b;
mem_array[37581] = 16'ha4c8;
mem_array[37580] = 16'h3cf1;
mem_array[37583] = 16'h87b6;
mem_array[37582] = 16'hbd80;
mem_array[37585] = 16'h29c8;
mem_array[37584] = 16'h3ebb;
mem_array[37587] = 16'h2bac;
mem_array[37586] = 16'h3eb0;
mem_array[37589] = 16'h3f94;
mem_array[37588] = 16'hbe35;
mem_array[37591] = 16'h3141;
mem_array[37590] = 16'hbe5f;
mem_array[37593] = 16'ha681;
mem_array[37592] = 16'hbec2;
mem_array[37595] = 16'hce4a;
mem_array[37594] = 16'hbe3d;
mem_array[37597] = 16'hdefb;
mem_array[37596] = 16'h3d99;
mem_array[37599] = 16'h95b6;
mem_array[37598] = 16'hbf01;
mem_array[37601] = 16'h84e3;
mem_array[37600] = 16'hbe50;
mem_array[37603] = 16'hd1d8;
mem_array[37602] = 16'hbbdd;
mem_array[37605] = 16'hcf42;
mem_array[37604] = 16'h3deb;
mem_array[37607] = 16'hbfc0;
mem_array[37606] = 16'hbe67;
mem_array[37609] = 16'h82d8;
mem_array[37608] = 16'h3b6b;
mem_array[37611] = 16'h8732;
mem_array[37610] = 16'h3e41;
mem_array[37613] = 16'had6b;
mem_array[37612] = 16'h3e01;
mem_array[37615] = 16'h793f;
mem_array[37614] = 16'h3d2e;
mem_array[37617] = 16'hdf9c;
mem_array[37616] = 16'hbd56;
mem_array[37619] = 16'h9311;
mem_array[37618] = 16'hbe57;
mem_array[37621] = 16'ha6e9;
mem_array[37620] = 16'hbeb3;
mem_array[37623] = 16'hc2fc;
mem_array[37622] = 16'hbe1e;
mem_array[37625] = 16'h37a5;
mem_array[37624] = 16'h3eae;
mem_array[37627] = 16'hc126;
mem_array[37626] = 16'h3e22;
mem_array[37629] = 16'h6316;
mem_array[37628] = 16'hbd7d;
mem_array[37631] = 16'h4982;
mem_array[37630] = 16'hbea4;
mem_array[37633] = 16'h44b9;
mem_array[37632] = 16'h3d36;
mem_array[37635] = 16'h22a9;
mem_array[37634] = 16'h3cd3;
mem_array[37637] = 16'h6f13;
mem_array[37636] = 16'hbe8b;
mem_array[37639] = 16'h473b;
mem_array[37638] = 16'hbeb9;
mem_array[37641] = 16'h6998;
mem_array[37640] = 16'hbd03;
mem_array[37643] = 16'h4056;
mem_array[37642] = 16'hbd48;
mem_array[37645] = 16'he4c3;
mem_array[37644] = 16'h3eb8;
mem_array[37647] = 16'h5f12;
mem_array[37646] = 16'h3e64;
mem_array[37649] = 16'h9ac6;
mem_array[37648] = 16'hbe2e;
mem_array[37651] = 16'hea52;
mem_array[37650] = 16'hbe64;
mem_array[37653] = 16'h986a;
mem_array[37652] = 16'hbbbd;
mem_array[37655] = 16'h588a;
mem_array[37654] = 16'h3cf9;
mem_array[37657] = 16'h83cf;
mem_array[37656] = 16'hbec1;
mem_array[37659] = 16'h26d0;
mem_array[37658] = 16'hbcf1;
mem_array[37661] = 16'h3c84;
mem_array[37660] = 16'hbe92;
mem_array[37663] = 16'h316d;
mem_array[37662] = 16'h3dce;
mem_array[37665] = 16'h7a8c;
mem_array[37664] = 16'hbe88;
mem_array[37667] = 16'had8f;
mem_array[37666] = 16'h3b99;
mem_array[37669] = 16'hbf7b;
mem_array[37668] = 16'hbd33;
mem_array[37671] = 16'h2acd;
mem_array[37670] = 16'h3d21;
mem_array[37673] = 16'h04c2;
mem_array[37672] = 16'h3e95;
mem_array[37675] = 16'ha3f4;
mem_array[37674] = 16'h3dc0;
mem_array[37677] = 16'h3be8;
mem_array[37676] = 16'hbcc2;
mem_array[37679] = 16'h5c5b;
mem_array[37678] = 16'hbd8a;
mem_array[37681] = 16'h97f2;
mem_array[37680] = 16'hbef3;
mem_array[37683] = 16'hfbd4;
mem_array[37682] = 16'hbd05;
mem_array[37685] = 16'h1aa6;
mem_array[37684] = 16'hbd39;
mem_array[37687] = 16'h1d03;
mem_array[37686] = 16'hbcea;
mem_array[37689] = 16'h5b03;
mem_array[37688] = 16'hbca6;
mem_array[37691] = 16'h680b;
mem_array[37690] = 16'hbdc6;
mem_array[37693] = 16'h38e4;
mem_array[37692] = 16'hbe3c;
mem_array[37695] = 16'haec2;
mem_array[37694] = 16'hbe38;
mem_array[37697] = 16'h1b90;
mem_array[37696] = 16'h3e24;
mem_array[37699] = 16'h2cb2;
mem_array[37698] = 16'hbd99;
mem_array[37701] = 16'hdbeb;
mem_array[37700] = 16'hbd8d;
mem_array[37703] = 16'he3ee;
mem_array[37702] = 16'hbce1;
mem_array[37705] = 16'h9830;
mem_array[37704] = 16'h3b21;
mem_array[37707] = 16'hf0b1;
mem_array[37706] = 16'h3d0e;
mem_array[37709] = 16'hc792;
mem_array[37708] = 16'hbe25;
mem_array[37711] = 16'h98c5;
mem_array[37710] = 16'hbd09;
mem_array[37713] = 16'h2503;
mem_array[37712] = 16'hbe8e;
mem_array[37715] = 16'hf609;
mem_array[37714] = 16'h3c81;
mem_array[37717] = 16'hcb87;
mem_array[37716] = 16'hbecb;
mem_array[37719] = 16'h4ab2;
mem_array[37718] = 16'h3bb4;
mem_array[37721] = 16'h97e7;
mem_array[37720] = 16'hbe9d;
mem_array[37723] = 16'hdaf7;
mem_array[37722] = 16'hbcac;
mem_array[37725] = 16'h7376;
mem_array[37724] = 16'h3e1a;
mem_array[37727] = 16'h4a43;
mem_array[37726] = 16'hbe07;
mem_array[37729] = 16'h4bcb;
mem_array[37728] = 16'hbe82;
mem_array[37731] = 16'h7278;
mem_array[37730] = 16'hbe5e;
mem_array[37733] = 16'hce40;
mem_array[37732] = 16'h3e4b;
mem_array[37735] = 16'h982a;
mem_array[37734] = 16'hbc92;
mem_array[37737] = 16'h193c;
mem_array[37736] = 16'h3e36;
mem_array[37739] = 16'h0e99;
mem_array[37738] = 16'h3e46;
mem_array[37741] = 16'h4723;
mem_array[37740] = 16'h3cd9;
mem_array[37743] = 16'h40e4;
mem_array[37742] = 16'hbd96;
mem_array[37745] = 16'h5f80;
mem_array[37744] = 16'h3e32;
mem_array[37747] = 16'h0fad;
mem_array[37746] = 16'h3cba;
mem_array[37749] = 16'h5936;
mem_array[37748] = 16'hbee0;
mem_array[37751] = 16'h45e0;
mem_array[37750] = 16'hbd8b;
mem_array[37753] = 16'h3b2b;
mem_array[37752] = 16'hbddc;
mem_array[37755] = 16'h1a59;
mem_array[37754] = 16'hbe80;
mem_array[37757] = 16'h1a83;
mem_array[37756] = 16'hbeb0;
mem_array[37759] = 16'hd840;
mem_array[37758] = 16'hbdde;
mem_array[37761] = 16'h8508;
mem_array[37760] = 16'h3c5d;
mem_array[37763] = 16'h1fab;
mem_array[37762] = 16'hbd82;
mem_array[37765] = 16'h474c;
mem_array[37764] = 16'hbe91;
mem_array[37767] = 16'ha563;
mem_array[37766] = 16'hbe76;
mem_array[37769] = 16'h4ce4;
mem_array[37768] = 16'hbe20;
mem_array[37771] = 16'h6f51;
mem_array[37770] = 16'hbe0c;
mem_array[37773] = 16'h0feb;
mem_array[37772] = 16'hbd96;
mem_array[37775] = 16'hb9f6;
mem_array[37774] = 16'hbd6c;
mem_array[37777] = 16'h9698;
mem_array[37776] = 16'hbea4;
mem_array[37779] = 16'h7ffe;
mem_array[37778] = 16'hbe5a;
mem_array[37781] = 16'h658c;
mem_array[37780] = 16'hbee6;
mem_array[37783] = 16'h1145;
mem_array[37782] = 16'hbd0b;
mem_array[37785] = 16'h4761;
mem_array[37784] = 16'h3e44;
mem_array[37787] = 16'h7902;
mem_array[37786] = 16'h3d27;
mem_array[37789] = 16'h544e;
mem_array[37788] = 16'hbccb;
mem_array[37791] = 16'h79e1;
mem_array[37790] = 16'h3d81;
mem_array[37793] = 16'h9f6a;
mem_array[37792] = 16'h3e3a;
mem_array[37795] = 16'h6002;
mem_array[37794] = 16'hbca7;
mem_array[37797] = 16'h0292;
mem_array[37796] = 16'hbece;
mem_array[37799] = 16'h2f88;
mem_array[37798] = 16'hbd40;
mem_array[37801] = 16'he2b4;
mem_array[37800] = 16'h3e65;
mem_array[37803] = 16'hee26;
mem_array[37802] = 16'h3e20;
mem_array[37805] = 16'h93aa;
mem_array[37804] = 16'h3dee;
mem_array[37807] = 16'h1f60;
mem_array[37806] = 16'h3d86;
mem_array[37809] = 16'hc430;
mem_array[37808] = 16'hbfdb;
mem_array[37811] = 16'hd461;
mem_array[37810] = 16'hbd10;
mem_array[37813] = 16'hb5f0;
mem_array[37812] = 16'hbdb3;
mem_array[37815] = 16'he122;
mem_array[37814] = 16'hbeb2;
mem_array[37817] = 16'hb765;
mem_array[37816] = 16'hbd8f;
mem_array[37819] = 16'h438e;
mem_array[37818] = 16'hbe29;
mem_array[37821] = 16'hd3d5;
mem_array[37820] = 16'h3ca7;
mem_array[37823] = 16'hd383;
mem_array[37822] = 16'h3c97;
mem_array[37825] = 16'hdafe;
mem_array[37824] = 16'hbeb2;
mem_array[37827] = 16'h25f5;
mem_array[37826] = 16'hbef3;
mem_array[37829] = 16'heaad;
mem_array[37828] = 16'hbec7;
mem_array[37831] = 16'hd12e;
mem_array[37830] = 16'hbe3f;
mem_array[37833] = 16'hd08c;
mem_array[37832] = 16'h3eed;
mem_array[37835] = 16'hbc72;
mem_array[37834] = 16'hbe0e;
mem_array[37837] = 16'h9f8f;
mem_array[37836] = 16'hbe9a;
mem_array[37839] = 16'h4ae6;
mem_array[37838] = 16'hbe34;
mem_array[37841] = 16'hb6c6;
mem_array[37840] = 16'hbe84;
mem_array[37843] = 16'h55a7;
mem_array[37842] = 16'hbd35;
mem_array[37845] = 16'h0f11;
mem_array[37844] = 16'hbd87;
mem_array[37847] = 16'h0cd8;
mem_array[37846] = 16'hba9f;
mem_array[37849] = 16'hd8db;
mem_array[37848] = 16'hbe4e;
mem_array[37851] = 16'h0892;
mem_array[37850] = 16'hbeb1;
mem_array[37853] = 16'hbe04;
mem_array[37852] = 16'h3df0;
mem_array[37855] = 16'ha584;
mem_array[37854] = 16'h3b86;
mem_array[37857] = 16'hc315;
mem_array[37856] = 16'hbf8f;
mem_array[37859] = 16'h3218;
mem_array[37858] = 16'h3bd4;
mem_array[37861] = 16'h1a7b;
mem_array[37860] = 16'hbf0d;
mem_array[37863] = 16'hc306;
mem_array[37862] = 16'h3da2;
mem_array[37865] = 16'h927e;
mem_array[37864] = 16'hbe10;
mem_array[37867] = 16'h4a48;
mem_array[37866] = 16'hbd7a;
mem_array[37869] = 16'haccd;
mem_array[37868] = 16'hbe14;
mem_array[37871] = 16'hf166;
mem_array[37870] = 16'hbe07;
mem_array[37873] = 16'h1c08;
mem_array[37872] = 16'h3d53;
mem_array[37875] = 16'h774b;
mem_array[37874] = 16'hbcb6;
mem_array[37877] = 16'ha4aa;
mem_array[37876] = 16'hbe9c;
mem_array[37879] = 16'h59bc;
mem_array[37878] = 16'h3c88;
mem_array[37881] = 16'h9bc3;
mem_array[37880] = 16'h3d59;
mem_array[37883] = 16'hee6e;
mem_array[37882] = 16'hbc5a;
mem_array[37885] = 16'h136d;
mem_array[37884] = 16'hbf09;
mem_array[37887] = 16'h62a8;
mem_array[37886] = 16'hbf02;
mem_array[37889] = 16'hde27;
mem_array[37888] = 16'h3d70;
mem_array[37891] = 16'h42d5;
mem_array[37890] = 16'hbe34;
mem_array[37893] = 16'h10fa;
mem_array[37892] = 16'h3e88;
mem_array[37895] = 16'h35cb;
mem_array[37894] = 16'hbc9c;
mem_array[37897] = 16'hc49e;
mem_array[37896] = 16'hbe72;
mem_array[37899] = 16'h87d6;
mem_array[37898] = 16'hbe2e;
mem_array[37901] = 16'hc1dd;
mem_array[37900] = 16'hbe00;
mem_array[37903] = 16'hde4e;
mem_array[37902] = 16'hbe2e;
mem_array[37905] = 16'h1dc1;
mem_array[37904] = 16'h3e29;
mem_array[37907] = 16'h87ff;
mem_array[37906] = 16'hbe10;
mem_array[37909] = 16'h690d;
mem_array[37908] = 16'h3dc9;
mem_array[37911] = 16'h0da1;
mem_array[37910] = 16'h3e58;
mem_array[37913] = 16'h0f24;
mem_array[37912] = 16'h3d79;
mem_array[37915] = 16'hcbc3;
mem_array[37914] = 16'hbe33;
mem_array[37917] = 16'h3d22;
mem_array[37916] = 16'hbf28;
mem_array[37919] = 16'h78dc;
mem_array[37918] = 16'h3e80;
mem_array[37921] = 16'h2e28;
mem_array[37920] = 16'h3e66;
mem_array[37923] = 16'h96ba;
mem_array[37922] = 16'h3cf2;
mem_array[37925] = 16'h6335;
mem_array[37924] = 16'hbead;
mem_array[37927] = 16'h09a4;
mem_array[37926] = 16'hbc23;
mem_array[37929] = 16'h2c31;
mem_array[37928] = 16'hbe9c;
mem_array[37931] = 16'h6654;
mem_array[37930] = 16'h3d13;
mem_array[37933] = 16'hc4e5;
mem_array[37932] = 16'h3db7;
mem_array[37935] = 16'hac23;
mem_array[37934] = 16'hbdb8;
mem_array[37937] = 16'hd6f9;
mem_array[37936] = 16'hbf5b;
mem_array[37939] = 16'hc799;
mem_array[37938] = 16'h3dfa;
mem_array[37941] = 16'h8e9d;
mem_array[37940] = 16'hbd5f;
mem_array[37943] = 16'h9d64;
mem_array[37942] = 16'hbdf9;
mem_array[37945] = 16'h52a4;
mem_array[37944] = 16'hbd5c;
mem_array[37947] = 16'h7787;
mem_array[37946] = 16'hbeec;
mem_array[37949] = 16'h25a0;
mem_array[37948] = 16'h3e07;
mem_array[37951] = 16'h2e05;
mem_array[37950] = 16'hbe4c;
mem_array[37953] = 16'h11f0;
mem_array[37952] = 16'h3ed4;
mem_array[37955] = 16'h5d56;
mem_array[37954] = 16'hbe4f;
mem_array[37957] = 16'h216f;
mem_array[37956] = 16'hbe80;
mem_array[37959] = 16'hb649;
mem_array[37958] = 16'hbed7;
mem_array[37961] = 16'hf576;
mem_array[37960] = 16'h3ed3;
mem_array[37963] = 16'hdb95;
mem_array[37962] = 16'h3c93;
mem_array[37965] = 16'h6a0c;
mem_array[37964] = 16'h3df4;
mem_array[37967] = 16'h30fb;
mem_array[37966] = 16'h3bf5;
mem_array[37969] = 16'ha971;
mem_array[37968] = 16'h3e21;
mem_array[37971] = 16'h47ab;
mem_array[37970] = 16'hbca6;
mem_array[37973] = 16'h8791;
mem_array[37972] = 16'hbd27;
mem_array[37975] = 16'hbce0;
mem_array[37974] = 16'hbe31;
mem_array[37977] = 16'h0ab1;
mem_array[37976] = 16'hbf24;
mem_array[37979] = 16'h10d7;
mem_array[37978] = 16'h3e65;
mem_array[37981] = 16'hf283;
mem_array[37980] = 16'hbefd;
mem_array[37983] = 16'h1929;
mem_array[37982] = 16'h3e9b;
mem_array[37985] = 16'hbcc0;
mem_array[37984] = 16'hbc25;
mem_array[37987] = 16'h1f8c;
mem_array[37986] = 16'h3e4d;
mem_array[37989] = 16'heacf;
mem_array[37988] = 16'hbea6;
mem_array[37991] = 16'ha7d0;
mem_array[37990] = 16'h3db6;
mem_array[37993] = 16'hc135;
mem_array[37992] = 16'hbe1d;
mem_array[37995] = 16'hbffb;
mem_array[37994] = 16'h3e94;
mem_array[37997] = 16'h1f20;
mem_array[37996] = 16'hbf5d;
mem_array[37999] = 16'h427b;
mem_array[37998] = 16'hbea1;
mem_array[38001] = 16'h66fb;
mem_array[38000] = 16'hbd38;
mem_array[38003] = 16'h19ef;
mem_array[38002] = 16'hbcf4;
mem_array[38005] = 16'h4338;
mem_array[38004] = 16'hbd95;
mem_array[38007] = 16'he774;
mem_array[38006] = 16'hbdb5;
mem_array[38009] = 16'h91f5;
mem_array[38008] = 16'h3ee2;
mem_array[38011] = 16'hdd5d;
mem_array[38010] = 16'hbe50;
mem_array[38013] = 16'h7668;
mem_array[38012] = 16'h3ecf;
mem_array[38015] = 16'hcf2c;
mem_array[38014] = 16'hbe1f;
mem_array[38017] = 16'h6e5d;
mem_array[38016] = 16'hbe65;
mem_array[38019] = 16'h99a8;
mem_array[38018] = 16'hbe37;
mem_array[38021] = 16'h4df6;
mem_array[38020] = 16'hbdea;
mem_array[38023] = 16'h64f1;
mem_array[38022] = 16'h3da6;
mem_array[38025] = 16'h8a57;
mem_array[38024] = 16'h3d2c;
mem_array[38027] = 16'h5406;
mem_array[38026] = 16'h3ddb;
mem_array[38029] = 16'h18fa;
mem_array[38028] = 16'h3dbe;
mem_array[38031] = 16'hf235;
mem_array[38030] = 16'h3e11;
mem_array[38033] = 16'ha91f;
mem_array[38032] = 16'h3d8f;
mem_array[38035] = 16'h48df;
mem_array[38034] = 16'hbd82;
mem_array[38037] = 16'he4ae;
mem_array[38036] = 16'hbf50;
mem_array[38039] = 16'he429;
mem_array[38038] = 16'hbe26;
mem_array[38041] = 16'hc064;
mem_array[38040] = 16'hbf7f;
mem_array[38043] = 16'h0042;
mem_array[38042] = 16'h3e8f;
mem_array[38045] = 16'h01a2;
mem_array[38044] = 16'hbd2a;
mem_array[38047] = 16'hf70d;
mem_array[38046] = 16'h3e89;
mem_array[38049] = 16'h425c;
mem_array[38048] = 16'h3f2c;
mem_array[38051] = 16'h2fdb;
mem_array[38050] = 16'h3e82;
mem_array[38053] = 16'hbb71;
mem_array[38052] = 16'h3dd6;
mem_array[38055] = 16'h2943;
mem_array[38054] = 16'hbe31;
mem_array[38057] = 16'haee9;
mem_array[38056] = 16'hbeb6;
mem_array[38059] = 16'ha877;
mem_array[38058] = 16'h3efc;
mem_array[38061] = 16'hd52e;
mem_array[38060] = 16'hbd6c;
mem_array[38063] = 16'h82f6;
mem_array[38062] = 16'hbdaa;
mem_array[38065] = 16'he279;
mem_array[38064] = 16'hbd1c;
mem_array[38067] = 16'hce30;
mem_array[38066] = 16'hbe1f;
mem_array[38069] = 16'h8172;
mem_array[38068] = 16'h3ec6;
mem_array[38071] = 16'h142e;
mem_array[38070] = 16'hbd52;
mem_array[38073] = 16'h2858;
mem_array[38072] = 16'h3f47;
mem_array[38075] = 16'h816f;
mem_array[38074] = 16'hbed7;
mem_array[38077] = 16'h6551;
mem_array[38076] = 16'hbe80;
mem_array[38079] = 16'h3659;
mem_array[38078] = 16'hbe01;
mem_array[38081] = 16'hf9d6;
mem_array[38080] = 16'hbe24;
mem_array[38083] = 16'hccf1;
mem_array[38082] = 16'hbdeb;
mem_array[38085] = 16'h1d67;
mem_array[38084] = 16'hbeef;
mem_array[38087] = 16'h6f1b;
mem_array[38086] = 16'hbe09;
mem_array[38089] = 16'h2ca1;
mem_array[38088] = 16'hbed5;
mem_array[38091] = 16'hae20;
mem_array[38090] = 16'hbeb9;
mem_array[38093] = 16'hf2cd;
mem_array[38092] = 16'h3e56;
mem_array[38095] = 16'hefe4;
mem_array[38094] = 16'h3e06;
mem_array[38097] = 16'h5a33;
mem_array[38096] = 16'hbeb0;
mem_array[38099] = 16'hb183;
mem_array[38098] = 16'hbd9e;
mem_array[38101] = 16'h0434;
mem_array[38100] = 16'hbe17;
mem_array[38103] = 16'hab3d;
mem_array[38102] = 16'h3e9a;
mem_array[38105] = 16'h4d4b;
mem_array[38104] = 16'h3eef;
mem_array[38107] = 16'h966f;
mem_array[38106] = 16'hbd4a;
mem_array[38109] = 16'hc71c;
mem_array[38108] = 16'h3e69;
mem_array[38111] = 16'h4c58;
mem_array[38110] = 16'h3e3c;
mem_array[38113] = 16'hea6d;
mem_array[38112] = 16'h3e63;
mem_array[38115] = 16'hcdf3;
mem_array[38114] = 16'hbed5;
mem_array[38117] = 16'h6bbf;
mem_array[38116] = 16'hbfab;
mem_array[38119] = 16'hbcc7;
mem_array[38118] = 16'hbe05;
mem_array[38121] = 16'ha759;
mem_array[38120] = 16'h3cd7;
mem_array[38123] = 16'ha951;
mem_array[38122] = 16'h3d01;
mem_array[38125] = 16'h29fc;
mem_array[38124] = 16'hbf0d;
mem_array[38127] = 16'ha373;
mem_array[38126] = 16'h3d95;
mem_array[38129] = 16'h14fa;
mem_array[38128] = 16'h3e1d;
mem_array[38131] = 16'hb103;
mem_array[38130] = 16'hbd9c;
mem_array[38133] = 16'ha91d;
mem_array[38132] = 16'h3efd;
mem_array[38135] = 16'heced;
mem_array[38134] = 16'hbd8d;
mem_array[38137] = 16'h0e82;
mem_array[38136] = 16'hbdca;
mem_array[38139] = 16'hc395;
mem_array[38138] = 16'hbe18;
mem_array[38141] = 16'haa3b;
mem_array[38140] = 16'h3f07;
mem_array[38143] = 16'h48bb;
mem_array[38142] = 16'hbefc;
mem_array[38145] = 16'hee76;
mem_array[38144] = 16'hbed8;
mem_array[38147] = 16'hd321;
mem_array[38146] = 16'hbe10;
mem_array[38149] = 16'h5a4a;
mem_array[38148] = 16'h3e82;
mem_array[38151] = 16'hab3e;
mem_array[38150] = 16'hbf3c;
mem_array[38153] = 16'hbca2;
mem_array[38152] = 16'h3ddf;
mem_array[38155] = 16'h292f;
mem_array[38154] = 16'hbe27;
mem_array[38157] = 16'hd722;
mem_array[38156] = 16'hbe4c;
mem_array[38159] = 16'ha652;
mem_array[38158] = 16'h3df3;
mem_array[38161] = 16'h0996;
mem_array[38160] = 16'hbee6;
mem_array[38163] = 16'h8e47;
mem_array[38162] = 16'h3e24;
mem_array[38165] = 16'h55f2;
mem_array[38164] = 16'hbc4b;
mem_array[38167] = 16'h8f7d;
mem_array[38166] = 16'h3ea7;
mem_array[38169] = 16'h9bae;
mem_array[38168] = 16'h3f09;
mem_array[38171] = 16'h391d;
mem_array[38170] = 16'h3e89;
mem_array[38173] = 16'he480;
mem_array[38172] = 16'h3d34;
mem_array[38175] = 16'he48b;
mem_array[38174] = 16'hbe32;
mem_array[38177] = 16'h4d3e;
mem_array[38176] = 16'hbf7b;
mem_array[38179] = 16'h5747;
mem_array[38178] = 16'hbd60;
mem_array[38181] = 16'hf740;
mem_array[38180] = 16'h3ca0;
mem_array[38183] = 16'h3006;
mem_array[38182] = 16'hbc4b;
mem_array[38185] = 16'hda72;
mem_array[38184] = 16'hbe43;
mem_array[38187] = 16'hc7f2;
mem_array[38186] = 16'h3df2;
mem_array[38189] = 16'h0ed1;
mem_array[38188] = 16'hbe04;
mem_array[38191] = 16'h2d97;
mem_array[38190] = 16'h3dc3;
mem_array[38193] = 16'h7d33;
mem_array[38192] = 16'hbeb9;
mem_array[38195] = 16'h1ef2;
mem_array[38194] = 16'hbe85;
mem_array[38197] = 16'h3372;
mem_array[38196] = 16'hbe55;
mem_array[38199] = 16'h5333;
mem_array[38198] = 16'hbe6b;
mem_array[38201] = 16'hc5db;
mem_array[38200] = 16'h3ead;
mem_array[38203] = 16'h56ac;
mem_array[38202] = 16'hbd5b;
mem_array[38205] = 16'h3699;
mem_array[38204] = 16'h3e44;
mem_array[38207] = 16'h6dc5;
mem_array[38206] = 16'hbe21;
mem_array[38209] = 16'hbd06;
mem_array[38208] = 16'h3da0;
mem_array[38211] = 16'hbf4a;
mem_array[38210] = 16'hbedf;
mem_array[38213] = 16'ha3ce;
mem_array[38212] = 16'h3e59;
mem_array[38215] = 16'h8ef1;
mem_array[38214] = 16'h3e2c;
mem_array[38217] = 16'hf2b0;
mem_array[38216] = 16'hbf05;
mem_array[38219] = 16'h1d53;
mem_array[38218] = 16'hbf0f;
mem_array[38221] = 16'ha6fa;
mem_array[38220] = 16'hbdb9;
mem_array[38223] = 16'hc0fe;
mem_array[38222] = 16'hbd77;
mem_array[38225] = 16'h2ecb;
mem_array[38224] = 16'h3ec8;
mem_array[38227] = 16'hb23e;
mem_array[38226] = 16'hbe87;
mem_array[38229] = 16'h6777;
mem_array[38228] = 16'h3eb7;
mem_array[38231] = 16'had97;
mem_array[38230] = 16'hbcbe;
mem_array[38233] = 16'h786f;
mem_array[38232] = 16'hbea9;
mem_array[38235] = 16'h7fba;
mem_array[38234] = 16'hbf81;
mem_array[38237] = 16'h7ee9;
mem_array[38236] = 16'hbf61;
mem_array[38239] = 16'h9556;
mem_array[38238] = 16'h3e33;
mem_array[38241] = 16'hd93d;
mem_array[38240] = 16'h3d66;
mem_array[38243] = 16'h9583;
mem_array[38242] = 16'h3ca6;
mem_array[38245] = 16'hed5f;
mem_array[38244] = 16'hbe2c;
mem_array[38247] = 16'h8559;
mem_array[38246] = 16'h3e40;
mem_array[38249] = 16'hf135;
mem_array[38248] = 16'h3ec1;
mem_array[38251] = 16'ha3f0;
mem_array[38250] = 16'h3c0f;
mem_array[38253] = 16'hea8e;
mem_array[38252] = 16'h3d4e;
mem_array[38255] = 16'h4bff;
mem_array[38254] = 16'hbdeb;
mem_array[38257] = 16'h899f;
mem_array[38256] = 16'hbee1;
mem_array[38259] = 16'hb765;
mem_array[38258] = 16'h3cfe;
mem_array[38261] = 16'hb05d;
mem_array[38260] = 16'h3db5;
mem_array[38263] = 16'ha513;
mem_array[38262] = 16'hbd4d;
mem_array[38265] = 16'ha57d;
mem_array[38264] = 16'hbf2e;
mem_array[38267] = 16'h368d;
mem_array[38266] = 16'h3e85;
mem_array[38269] = 16'hbfda;
mem_array[38268] = 16'hbe82;
mem_array[38271] = 16'h36dc;
mem_array[38270] = 16'hbe7f;
mem_array[38273] = 16'h47d8;
mem_array[38272] = 16'hbd9e;
mem_array[38275] = 16'h620c;
mem_array[38274] = 16'h3e20;
mem_array[38277] = 16'h208d;
mem_array[38276] = 16'hbf25;
mem_array[38279] = 16'habf7;
mem_array[38278] = 16'hbda3;
mem_array[38281] = 16'h653a;
mem_array[38280] = 16'h3ebe;
mem_array[38283] = 16'h440f;
mem_array[38282] = 16'hbe94;
mem_array[38285] = 16'h4d5b;
mem_array[38284] = 16'h3e79;
mem_array[38287] = 16'h712c;
mem_array[38286] = 16'h3d51;
mem_array[38289] = 16'hae1c;
mem_array[38288] = 16'h3d80;
mem_array[38291] = 16'h4d28;
mem_array[38290] = 16'hbf12;
mem_array[38293] = 16'ha955;
mem_array[38292] = 16'h3cb6;
mem_array[38295] = 16'hed1a;
mem_array[38294] = 16'hbf84;
mem_array[38297] = 16'hb0c6;
mem_array[38296] = 16'hbf57;
mem_array[38299] = 16'he57e;
mem_array[38298] = 16'h3d37;
mem_array[38301] = 16'hfc02;
mem_array[38300] = 16'h3ba5;
mem_array[38303] = 16'hc01d;
mem_array[38302] = 16'h3d10;
mem_array[38305] = 16'h3be4;
mem_array[38304] = 16'hbd92;
mem_array[38307] = 16'hf8d9;
mem_array[38306] = 16'h3ed2;
mem_array[38309] = 16'hd952;
mem_array[38308] = 16'h3e04;
mem_array[38311] = 16'hd7d3;
mem_array[38310] = 16'hbe7c;
mem_array[38313] = 16'h34ac;
mem_array[38312] = 16'h3e90;
mem_array[38315] = 16'h01e0;
mem_array[38314] = 16'h3dce;
mem_array[38317] = 16'h0fab;
mem_array[38316] = 16'hbe50;
mem_array[38319] = 16'h2f8f;
mem_array[38318] = 16'h3e46;
mem_array[38321] = 16'h4d99;
mem_array[38320] = 16'hbe77;
mem_array[38323] = 16'h1392;
mem_array[38322] = 16'h3e05;
mem_array[38325] = 16'h6a83;
mem_array[38324] = 16'hbe6b;
mem_array[38327] = 16'hcce0;
mem_array[38326] = 16'hbef6;
mem_array[38329] = 16'h05dd;
mem_array[38328] = 16'h3b44;
mem_array[38331] = 16'hd83e;
mem_array[38330] = 16'hbef8;
mem_array[38333] = 16'h275d;
mem_array[38332] = 16'h3ef5;
mem_array[38335] = 16'he12f;
mem_array[38334] = 16'h3e44;
mem_array[38337] = 16'heffc;
mem_array[38336] = 16'hbdc6;
mem_array[38339] = 16'hbca2;
mem_array[38338] = 16'hbdaa;
mem_array[38341] = 16'h40ed;
mem_array[38340] = 16'h3edf;
mem_array[38343] = 16'h8c9c;
mem_array[38342] = 16'h3d13;
mem_array[38345] = 16'h24d4;
mem_array[38344] = 16'h3e2e;
mem_array[38347] = 16'h6d93;
mem_array[38346] = 16'hbf15;
mem_array[38349] = 16'hdfc3;
mem_array[38348] = 16'h3eb7;
mem_array[38351] = 16'h02d3;
mem_array[38350] = 16'hbe98;
mem_array[38353] = 16'h672c;
mem_array[38352] = 16'h3f57;
mem_array[38355] = 16'h6b4a;
mem_array[38354] = 16'h3edb;
mem_array[38357] = 16'h0fc3;
mem_array[38356] = 16'h3db4;
mem_array[38359] = 16'h918e;
mem_array[38358] = 16'h3f01;
mem_array[38361] = 16'h8ae2;
mem_array[38360] = 16'h3d1a;
mem_array[38363] = 16'hcded;
mem_array[38362] = 16'h3c19;
mem_array[38365] = 16'hb554;
mem_array[38364] = 16'hbf89;
mem_array[38367] = 16'h5b8f;
mem_array[38366] = 16'hbdcb;
mem_array[38369] = 16'ha02e;
mem_array[38368] = 16'hbd54;
mem_array[38371] = 16'h0b2c;
mem_array[38370] = 16'hbd00;
mem_array[38373] = 16'hf578;
mem_array[38372] = 16'hbedf;
mem_array[38375] = 16'h47aa;
mem_array[38374] = 16'hbf3c;
mem_array[38377] = 16'h312d;
mem_array[38376] = 16'hbd8a;
mem_array[38379] = 16'h121a;
mem_array[38378] = 16'h3d05;
mem_array[38381] = 16'hd8be;
mem_array[38380] = 16'hbf70;
mem_array[38383] = 16'h08ec;
mem_array[38382] = 16'h3e65;
mem_array[38385] = 16'hf2aa;
mem_array[38384] = 16'hbe3a;
mem_array[38387] = 16'h50c6;
mem_array[38386] = 16'hbe7b;
mem_array[38389] = 16'h739f;
mem_array[38388] = 16'h3e8a;
mem_array[38391] = 16'h8b08;
mem_array[38390] = 16'hbf53;
mem_array[38393] = 16'hb647;
mem_array[38392] = 16'h3f81;
mem_array[38395] = 16'he479;
mem_array[38394] = 16'h3df5;
mem_array[38397] = 16'h72e7;
mem_array[38396] = 16'hbdaf;
mem_array[38399] = 16'hcf59;
mem_array[38398] = 16'hbf97;
mem_array[38401] = 16'h3621;
mem_array[38400] = 16'h3ee9;
mem_array[38403] = 16'hbc67;
mem_array[38402] = 16'hbcd1;
mem_array[38405] = 16'h4701;
mem_array[38404] = 16'h3e56;
mem_array[38407] = 16'hb237;
mem_array[38406] = 16'hbf5f;
mem_array[38409] = 16'h873e;
mem_array[38408] = 16'hbdef;
mem_array[38411] = 16'h6945;
mem_array[38410] = 16'hbf08;
mem_array[38413] = 16'h52fb;
mem_array[38412] = 16'hbe86;
mem_array[38415] = 16'hf727;
mem_array[38414] = 16'hbf2f;
mem_array[38417] = 16'h3ac5;
mem_array[38416] = 16'hbd6e;
mem_array[38419] = 16'he2f5;
mem_array[38418] = 16'h3f44;
mem_array[38421] = 16'h9359;
mem_array[38420] = 16'h3d66;
mem_array[38423] = 16'hd60d;
mem_array[38422] = 16'hbc80;
mem_array[38425] = 16'h3338;
mem_array[38424] = 16'hbf48;
mem_array[38427] = 16'h226b;
mem_array[38426] = 16'h3ee6;
mem_array[38429] = 16'h0f4d;
mem_array[38428] = 16'h3ef4;
mem_array[38431] = 16'h2f3a;
mem_array[38430] = 16'h3df3;
mem_array[38433] = 16'hb6e6;
mem_array[38432] = 16'h3f67;
mem_array[38435] = 16'hb400;
mem_array[38434] = 16'hbe9f;
mem_array[38437] = 16'h6062;
mem_array[38436] = 16'h3daf;
mem_array[38439] = 16'h900e;
mem_array[38438] = 16'hbe10;
mem_array[38441] = 16'h02c1;
mem_array[38440] = 16'hbf45;
mem_array[38443] = 16'hc5c1;
mem_array[38442] = 16'h3e30;
mem_array[38445] = 16'hc072;
mem_array[38444] = 16'hbf4f;
mem_array[38447] = 16'h19e4;
mem_array[38446] = 16'h3f54;
mem_array[38449] = 16'h9cf1;
mem_array[38448] = 16'hbe2b;
mem_array[38451] = 16'h8e14;
mem_array[38450] = 16'hbc3e;
mem_array[38453] = 16'h4dd1;
mem_array[38452] = 16'h3efc;
mem_array[38455] = 16'he526;
mem_array[38454] = 16'hbec1;
mem_array[38457] = 16'hfb86;
mem_array[38456] = 16'h3ec5;
mem_array[38459] = 16'h0fbb;
mem_array[38458] = 16'hbeb2;
mem_array[38461] = 16'h9eef;
mem_array[38460] = 16'h3cf1;
mem_array[38463] = 16'h95d3;
mem_array[38462] = 16'hbd45;
mem_array[38465] = 16'hbf13;
mem_array[38464] = 16'h3f48;
mem_array[38467] = 16'h83b8;
mem_array[38466] = 16'h3e10;
mem_array[38469] = 16'h0805;
mem_array[38468] = 16'hbe39;
mem_array[38471] = 16'hba9b;
mem_array[38470] = 16'hbe00;
mem_array[38473] = 16'h7c8b;
mem_array[38472] = 16'hbde2;
mem_array[38475] = 16'hd5e4;
mem_array[38474] = 16'hbe73;
mem_array[38477] = 16'hf270;
mem_array[38476] = 16'h3f08;
mem_array[38479] = 16'h33be;
mem_array[38478] = 16'h3fa3;
mem_array[38481] = 16'h3ebe;
mem_array[38480] = 16'hbd9b;
mem_array[38483] = 16'hc629;
mem_array[38482] = 16'h3d90;
mem_array[38485] = 16'h922e;
mem_array[38484] = 16'h3f3c;
mem_array[38487] = 16'hcac9;
mem_array[38486] = 16'hbf06;
mem_array[38489] = 16'h7e59;
mem_array[38488] = 16'h3ecb;
mem_array[38491] = 16'h6e58;
mem_array[38490] = 16'hbe77;
mem_array[38493] = 16'h7ce5;
mem_array[38492] = 16'h3fcb;
mem_array[38495] = 16'h83ec;
mem_array[38494] = 16'h3e05;
mem_array[38497] = 16'h3148;
mem_array[38496] = 16'h39aa;
mem_array[38499] = 16'h8d69;
mem_array[38498] = 16'hbe4f;
mem_array[38501] = 16'h280e;
mem_array[38500] = 16'hbf11;
mem_array[38503] = 16'hb106;
mem_array[38502] = 16'h3c9e;
mem_array[38505] = 16'hf825;
mem_array[38504] = 16'hbf27;
mem_array[38507] = 16'h1ad4;
mem_array[38506] = 16'h3f69;
mem_array[38509] = 16'hd1b0;
mem_array[38508] = 16'hbd86;
mem_array[38511] = 16'h2e79;
mem_array[38510] = 16'h3ec5;
mem_array[38513] = 16'hd45a;
mem_array[38512] = 16'h3e57;
mem_array[38515] = 16'h13f6;
mem_array[38514] = 16'hbf3c;
mem_array[38517] = 16'hedfa;
mem_array[38516] = 16'h3f2b;
mem_array[38519] = 16'hd1bd;
mem_array[38518] = 16'hbeb6;
mem_array[38521] = 16'h2ff6;
mem_array[38520] = 16'h3f54;
mem_array[38523] = 16'ha3cd;
mem_array[38522] = 16'h3dde;
mem_array[38525] = 16'he7e4;
mem_array[38524] = 16'h3ded;
mem_array[38527] = 16'h2dac;
mem_array[38526] = 16'h3fec;
mem_array[38529] = 16'h2a0a;
mem_array[38528] = 16'h3d49;
mem_array[38531] = 16'h67e7;
mem_array[38530] = 16'h3e5c;
mem_array[38533] = 16'h0d25;
mem_array[38532] = 16'hbeff;
mem_array[38535] = 16'hbcfb;
mem_array[38534] = 16'h3d8a;
mem_array[38537] = 16'h0a01;
mem_array[38536] = 16'hbd81;
mem_array[38539] = 16'ha387;
mem_array[38538] = 16'h3f79;
mem_array[38541] = 16'h96b0;
mem_array[38540] = 16'h3d14;
mem_array[38543] = 16'h2022;
mem_array[38542] = 16'hbda9;
mem_array[38545] = 16'hc61f;
mem_array[38544] = 16'h3fb3;
mem_array[38547] = 16'h219e;
mem_array[38546] = 16'hbfa2;
mem_array[38549] = 16'h6725;
mem_array[38548] = 16'h3c10;
mem_array[38551] = 16'h2efb;
mem_array[38550] = 16'hbf7c;
mem_array[38553] = 16'hd3b7;
mem_array[38552] = 16'h3eac;
mem_array[38555] = 16'h9f6c;
mem_array[38554] = 16'h3f4a;
mem_array[38557] = 16'h61ae;
mem_array[38556] = 16'hbf96;
mem_array[38559] = 16'h31bc;
mem_array[38558] = 16'h3ed2;
mem_array[38561] = 16'hbc22;
mem_array[38560] = 16'h3f26;
mem_array[38563] = 16'h3157;
mem_array[38562] = 16'h3ed3;
mem_array[38565] = 16'h6e23;
mem_array[38564] = 16'hbe25;
mem_array[38567] = 16'h2b01;
mem_array[38566] = 16'h3f5d;
mem_array[38569] = 16'hcf30;
mem_array[38568] = 16'h3e45;
mem_array[38571] = 16'h92ed;
mem_array[38570] = 16'h3d8d;
mem_array[38573] = 16'hfe8a;
mem_array[38572] = 16'hbf2c;
mem_array[38575] = 16'h2d24;
mem_array[38574] = 16'h3d93;
mem_array[38577] = 16'h09d6;
mem_array[38576] = 16'hbf24;
mem_array[38579] = 16'hf8e8;
mem_array[38578] = 16'h3f67;
mem_array[38581] = 16'hfcd4;
mem_array[38580] = 16'h3bb9;
mem_array[38583] = 16'hacc4;
mem_array[38582] = 16'hbbd8;
mem_array[38585] = 16'h5d52;
mem_array[38584] = 16'h3c28;
mem_array[38587] = 16'h856a;
mem_array[38586] = 16'hbd27;
mem_array[38589] = 16'hbda2;
mem_array[38588] = 16'hbc9b;
mem_array[38591] = 16'h344e;
mem_array[38590] = 16'hbbfe;
mem_array[38593] = 16'hf267;
mem_array[38592] = 16'h3da1;
mem_array[38595] = 16'he1e6;
mem_array[38594] = 16'h3c89;
mem_array[38597] = 16'h136c;
mem_array[38596] = 16'hbdba;
mem_array[38599] = 16'h7294;
mem_array[38598] = 16'hbcdb;
mem_array[38601] = 16'h56e2;
mem_array[38600] = 16'h3dae;
mem_array[38603] = 16'hbe11;
mem_array[38602] = 16'hbd31;
mem_array[38605] = 16'h12da;
mem_array[38604] = 16'h3dc3;
mem_array[38607] = 16'h66d9;
mem_array[38606] = 16'h3cf6;
mem_array[38609] = 16'h5c6a;
mem_array[38608] = 16'hbd6d;
mem_array[38611] = 16'h8165;
mem_array[38610] = 16'hbd84;
mem_array[38613] = 16'h6f3a;
mem_array[38612] = 16'h3d15;
mem_array[38615] = 16'h2feb;
mem_array[38614] = 16'h3cdf;
mem_array[38617] = 16'hac9e;
mem_array[38616] = 16'h3d4a;
mem_array[38619] = 16'h9885;
mem_array[38618] = 16'h3ddd;
mem_array[38621] = 16'hb4a4;
mem_array[38620] = 16'h3cef;
mem_array[38623] = 16'hf5d0;
mem_array[38622] = 16'hbdf7;
mem_array[38625] = 16'hfd56;
mem_array[38624] = 16'hbb86;
mem_array[38627] = 16'h64ca;
mem_array[38626] = 16'hbd9a;
mem_array[38629] = 16'h0a16;
mem_array[38628] = 16'h3d6e;
mem_array[38631] = 16'h1e13;
mem_array[38630] = 16'h3ccf;
mem_array[38633] = 16'h0ba3;
mem_array[38632] = 16'h3cdd;
mem_array[38635] = 16'h546d;
mem_array[38634] = 16'h3d8a;
mem_array[38637] = 16'he9b1;
mem_array[38636] = 16'hbd08;
mem_array[38639] = 16'he574;
mem_array[38638] = 16'hbcc5;
mem_array[38641] = 16'h36a5;
mem_array[38640] = 16'h3ceb;
mem_array[38643] = 16'h6712;
mem_array[38642] = 16'h3d8e;
mem_array[38645] = 16'h4715;
mem_array[38644] = 16'hbd96;
mem_array[38647] = 16'hf309;
mem_array[38646] = 16'h3d4e;
mem_array[38649] = 16'h1c13;
mem_array[38648] = 16'hbd46;
mem_array[38651] = 16'h5530;
mem_array[38650] = 16'h3d99;
mem_array[38653] = 16'h0fba;
mem_array[38652] = 16'h3cab;
mem_array[38655] = 16'h93ea;
mem_array[38654] = 16'hbd45;
mem_array[38657] = 16'h548e;
mem_array[38656] = 16'h3dbb;
mem_array[38659] = 16'h177c;
mem_array[38658] = 16'hbd68;
mem_array[38661] = 16'h0801;
mem_array[38660] = 16'h3d9a;
mem_array[38663] = 16'h1297;
mem_array[38662] = 16'h3bd1;
mem_array[38665] = 16'h4228;
mem_array[38664] = 16'hbc98;
mem_array[38667] = 16'h0978;
mem_array[38666] = 16'hbd04;
mem_array[38669] = 16'h0cee;
mem_array[38668] = 16'h3c4c;
mem_array[38671] = 16'h6708;
mem_array[38670] = 16'hbc01;
mem_array[38673] = 16'hd164;
mem_array[38672] = 16'hbcd4;
mem_array[38675] = 16'h3565;
mem_array[38674] = 16'h3d04;
mem_array[38677] = 16'h09d5;
mem_array[38676] = 16'h3caa;
mem_array[38679] = 16'h7822;
mem_array[38678] = 16'hbd3d;
mem_array[38681] = 16'h0a77;
mem_array[38680] = 16'h3cbb;
mem_array[38683] = 16'he208;
mem_array[38682] = 16'h3cf7;
mem_array[38685] = 16'h9cc5;
mem_array[38684] = 16'h3d84;
mem_array[38687] = 16'h3f78;
mem_array[38686] = 16'h3c8b;
mem_array[38689] = 16'hf870;
mem_array[38688] = 16'hbd8c;
mem_array[38691] = 16'h8d14;
mem_array[38690] = 16'hbdb4;
mem_array[38693] = 16'h0c84;
mem_array[38692] = 16'h3b84;
mem_array[38695] = 16'h97ab;
mem_array[38694] = 16'h3c24;
mem_array[38697] = 16'h06fd;
mem_array[38696] = 16'h3d7e;
mem_array[38699] = 16'h4faa;
mem_array[38698] = 16'hbdea;
mem_array[38701] = 16'hf14c;
mem_array[38700] = 16'h3c8a;
mem_array[38703] = 16'h8b72;
mem_array[38702] = 16'h3ca0;
mem_array[38705] = 16'h70ca;
mem_array[38704] = 16'hbc8b;
mem_array[38707] = 16'h55c7;
mem_array[38706] = 16'hbd42;
mem_array[38709] = 16'h7600;
mem_array[38708] = 16'hbd58;
mem_array[38711] = 16'h2a71;
mem_array[38710] = 16'hbd2f;
mem_array[38713] = 16'ha209;
mem_array[38712] = 16'hbdc5;
mem_array[38715] = 16'heabf;
mem_array[38714] = 16'hbd3e;
mem_array[38717] = 16'h9444;
mem_array[38716] = 16'h3cee;
mem_array[38719] = 16'hcc6b;
mem_array[38718] = 16'hbdde;
mem_array[38721] = 16'ha876;
mem_array[38720] = 16'h3d44;
mem_array[38723] = 16'hf00c;
mem_array[38722] = 16'h3cb7;
mem_array[38725] = 16'hab59;
mem_array[38724] = 16'hbab8;
mem_array[38727] = 16'had03;
mem_array[38726] = 16'hbd90;
mem_array[38729] = 16'hfff1;
mem_array[38728] = 16'h3bdb;
mem_array[38731] = 16'hd622;
mem_array[38730] = 16'h3cb5;
mem_array[38733] = 16'hec5d;
mem_array[38732] = 16'h3cb5;
mem_array[38735] = 16'h6dc8;
mem_array[38734] = 16'h3d45;
mem_array[38737] = 16'hd1d7;
mem_array[38736] = 16'h3d91;
mem_array[38739] = 16'hb704;
mem_array[38738] = 16'hbd81;
mem_array[38741] = 16'h3d1f;
mem_array[38740] = 16'hbd8b;
mem_array[38743] = 16'hb9f6;
mem_array[38742] = 16'hbd16;
mem_array[38745] = 16'hf5b1;
mem_array[38744] = 16'hbb4b;
mem_array[38747] = 16'h1f11;
mem_array[38746] = 16'hbd7c;
mem_array[38749] = 16'hd0fc;
mem_array[38748] = 16'h3c42;
mem_array[38751] = 16'h2d00;
mem_array[38750] = 16'hbcf2;
mem_array[38753] = 16'h578f;
mem_array[38752] = 16'h3d62;
mem_array[38755] = 16'hd5c1;
mem_array[38754] = 16'hbd34;
mem_array[38757] = 16'h818f;
mem_array[38756] = 16'h3ca5;
mem_array[38759] = 16'hccff;
mem_array[38758] = 16'h3d48;
mem_array[38761] = 16'h5229;
mem_array[38760] = 16'hbe14;
mem_array[38763] = 16'h68e1;
mem_array[38762] = 16'h3ec9;
mem_array[38765] = 16'h2bcf;
mem_array[38764] = 16'h3f20;
mem_array[38767] = 16'h35e3;
mem_array[38766] = 16'hbe08;
mem_array[38769] = 16'h4c7f;
mem_array[38768] = 16'hbec1;
mem_array[38771] = 16'h4568;
mem_array[38770] = 16'hbe86;
mem_array[38773] = 16'he0d9;
mem_array[38772] = 16'h3eb9;
mem_array[38775] = 16'h3bfd;
mem_array[38774] = 16'hbee0;
mem_array[38777] = 16'h5739;
mem_array[38776] = 16'h3e3c;
mem_array[38779] = 16'hbe96;
mem_array[38778] = 16'hbd32;
mem_array[38781] = 16'hb6c0;
mem_array[38780] = 16'h3d81;
mem_array[38783] = 16'h1992;
mem_array[38782] = 16'hbd05;
mem_array[38785] = 16'h0567;
mem_array[38784] = 16'hbecb;
mem_array[38787] = 16'h8a63;
mem_array[38786] = 16'h3f1c;
mem_array[38789] = 16'hf528;
mem_array[38788] = 16'h3eb2;
mem_array[38791] = 16'h5e4b;
mem_array[38790] = 16'hbe4c;
mem_array[38793] = 16'h6552;
mem_array[38792] = 16'h3bc9;
mem_array[38795] = 16'hf380;
mem_array[38794] = 16'h3d40;
mem_array[38797] = 16'h5912;
mem_array[38796] = 16'h3c84;
mem_array[38799] = 16'hdf02;
mem_array[38798] = 16'hbd30;
mem_array[38801] = 16'h95ca;
mem_array[38800] = 16'hbe71;
mem_array[38803] = 16'h8d68;
mem_array[38802] = 16'h3ca5;
mem_array[38805] = 16'hd1fe;
mem_array[38804] = 16'hbdc8;
mem_array[38807] = 16'h62ca;
mem_array[38806] = 16'hbf02;
mem_array[38809] = 16'hde12;
mem_array[38808] = 16'h3ee3;
mem_array[38811] = 16'h2196;
mem_array[38810] = 16'hbdd0;
mem_array[38813] = 16'h15bb;
mem_array[38812] = 16'h3f34;
mem_array[38815] = 16'h1fff;
mem_array[38814] = 16'h3f3d;
mem_array[38817] = 16'h1c51;
mem_array[38816] = 16'hbea8;
mem_array[38819] = 16'h5cae;
mem_array[38818] = 16'hbe66;
mem_array[38821] = 16'hc210;
mem_array[38820] = 16'hbf7b;
mem_array[38823] = 16'h08dd;
mem_array[38822] = 16'h3eb2;
mem_array[38825] = 16'h3552;
mem_array[38824] = 16'hbeab;
mem_array[38827] = 16'h68b6;
mem_array[38826] = 16'hbf48;
mem_array[38829] = 16'h9a95;
mem_array[38828] = 16'hbe87;
mem_array[38831] = 16'ha2d6;
mem_array[38830] = 16'hbf55;
mem_array[38833] = 16'hc44a;
mem_array[38832] = 16'h3ee7;
mem_array[38835] = 16'h437e;
mem_array[38834] = 16'hbe8e;
mem_array[38837] = 16'hf276;
mem_array[38836] = 16'hbe8e;
mem_array[38839] = 16'h3d09;
mem_array[38838] = 16'hbc7b;
mem_array[38841] = 16'ha17e;
mem_array[38840] = 16'h3d71;
mem_array[38843] = 16'h5b0d;
mem_array[38842] = 16'hbddb;
mem_array[38845] = 16'h13dd;
mem_array[38844] = 16'hbf51;
mem_array[38847] = 16'h7469;
mem_array[38846] = 16'hbf20;
mem_array[38849] = 16'he2d5;
mem_array[38848] = 16'hbe7f;
mem_array[38851] = 16'h7489;
mem_array[38850] = 16'hbe82;
mem_array[38853] = 16'hcd06;
mem_array[38852] = 16'h3f9e;
mem_array[38855] = 16'h3db1;
mem_array[38854] = 16'hbf37;
mem_array[38857] = 16'h4e6e;
mem_array[38856] = 16'h3c95;
mem_array[38859] = 16'hb271;
mem_array[38858] = 16'hbed7;
mem_array[38861] = 16'h857e;
mem_array[38860] = 16'hbf0e;
mem_array[38863] = 16'h6535;
mem_array[38862] = 16'h3e8e;
mem_array[38865] = 16'hdc9e;
mem_array[38864] = 16'hbdc1;
mem_array[38867] = 16'h42d7;
mem_array[38866] = 16'h3e29;
mem_array[38869] = 16'h3436;
mem_array[38868] = 16'hbea2;
mem_array[38871] = 16'hfded;
mem_array[38870] = 16'hbf54;
mem_array[38873] = 16'hc03a;
mem_array[38872] = 16'h3ed0;
mem_array[38875] = 16'h86a0;
mem_array[38874] = 16'hbd7b;
mem_array[38877] = 16'h8da2;
mem_array[38876] = 16'h3eb7;
mem_array[38879] = 16'h40e6;
mem_array[38878] = 16'h3e7f;
mem_array[38881] = 16'hccf7;
mem_array[38880] = 16'h3e2f;
mem_array[38883] = 16'hd08f;
mem_array[38882] = 16'h3f0d;
mem_array[38885] = 16'h748f;
mem_array[38884] = 16'hbf04;
mem_array[38887] = 16'ha79f;
mem_array[38886] = 16'hbf96;
mem_array[38889] = 16'hbba8;
mem_array[38888] = 16'hbd65;
mem_array[38891] = 16'hf690;
mem_array[38890] = 16'hbf19;
mem_array[38893] = 16'hfed2;
mem_array[38892] = 16'h3e8d;
mem_array[38895] = 16'h888e;
mem_array[38894] = 16'h3e50;
mem_array[38897] = 16'h5f74;
mem_array[38896] = 16'hbd82;
mem_array[38899] = 16'hbefb;
mem_array[38898] = 16'hbf36;
mem_array[38901] = 16'hb1d9;
mem_array[38900] = 16'hbb7a;
mem_array[38903] = 16'habb9;
mem_array[38902] = 16'hbc86;
mem_array[38905] = 16'h6d57;
mem_array[38904] = 16'hbf50;
mem_array[38907] = 16'he8a5;
mem_array[38906] = 16'hbe33;
mem_array[38909] = 16'hb0fc;
mem_array[38908] = 16'hbe35;
mem_array[38911] = 16'h0805;
mem_array[38910] = 16'hbd16;
mem_array[38913] = 16'h43e9;
mem_array[38912] = 16'h3e21;
mem_array[38915] = 16'h3aad;
mem_array[38914] = 16'hbf45;
mem_array[38917] = 16'h38d0;
mem_array[38916] = 16'hbfa7;
mem_array[38919] = 16'h6484;
mem_array[38918] = 16'hbf88;
mem_array[38921] = 16'h5c57;
mem_array[38920] = 16'hbfa8;
mem_array[38923] = 16'h2679;
mem_array[38922] = 16'h3f25;
mem_array[38925] = 16'h8a94;
mem_array[38924] = 16'hbcbf;
mem_array[38927] = 16'h8eb4;
mem_array[38926] = 16'h3ef8;
mem_array[38929] = 16'hf4ae;
mem_array[38928] = 16'h3f14;
mem_array[38931] = 16'hac9f;
mem_array[38930] = 16'hbd8f;
mem_array[38933] = 16'ha68b;
mem_array[38932] = 16'h3f47;
mem_array[38935] = 16'h4cb4;
mem_array[38934] = 16'h3f44;
mem_array[38937] = 16'hb2ab;
mem_array[38936] = 16'h3cc5;
mem_array[38939] = 16'haa96;
mem_array[38938] = 16'hbe92;
mem_array[38941] = 16'hb12f;
mem_array[38940] = 16'h3f0e;
mem_array[38943] = 16'h359e;
mem_array[38942] = 16'h3ed4;
mem_array[38945] = 16'h8290;
mem_array[38944] = 16'h3ded;
mem_array[38947] = 16'h345f;
mem_array[38946] = 16'h3ed1;
mem_array[38949] = 16'h9b49;
mem_array[38948] = 16'hbe29;
mem_array[38951] = 16'h8dd9;
mem_array[38950] = 16'h3f1e;
mem_array[38953] = 16'h3e9e;
mem_array[38952] = 16'h3e80;
mem_array[38955] = 16'h49b7;
mem_array[38954] = 16'h3d2d;
mem_array[38957] = 16'h2697;
mem_array[38956] = 16'h3d8a;
mem_array[38959] = 16'h7e12;
mem_array[38958] = 16'hbf71;
mem_array[38961] = 16'h86cb;
mem_array[38960] = 16'hbd28;
mem_array[38963] = 16'h0d02;
mem_array[38962] = 16'hbcf7;
mem_array[38965] = 16'h3221;
mem_array[38964] = 16'hbdbb;
mem_array[38967] = 16'h00ca;
mem_array[38966] = 16'h3eb8;
mem_array[38969] = 16'h776e;
mem_array[38968] = 16'h3eaa;
mem_array[38971] = 16'hc52b;
mem_array[38970] = 16'hbdc3;
mem_array[38973] = 16'h678a;
mem_array[38972] = 16'h3d80;
mem_array[38975] = 16'hcb8f;
mem_array[38974] = 16'hbf13;
mem_array[38977] = 16'h63b8;
mem_array[38976] = 16'hbf25;
mem_array[38979] = 16'h8cc0;
mem_array[38978] = 16'hbf03;
mem_array[38981] = 16'h0745;
mem_array[38980] = 16'hbf49;
mem_array[38983] = 16'h477c;
mem_array[38982] = 16'hbdde;
mem_array[38985] = 16'hde05;
mem_array[38984] = 16'hbead;
mem_array[38987] = 16'h728a;
mem_array[38986] = 16'hbee7;
mem_array[38989] = 16'h28b8;
mem_array[38988] = 16'h3f31;
mem_array[38991] = 16'h5da3;
mem_array[38990] = 16'h3f80;
mem_array[38993] = 16'h639e;
mem_array[38992] = 16'h3f59;
mem_array[38995] = 16'hdaae;
mem_array[38994] = 16'h3eff;
mem_array[38997] = 16'h5a54;
mem_array[38996] = 16'hbb16;
mem_array[38999] = 16'h3031;
mem_array[38998] = 16'hbee8;
mem_array[39001] = 16'ha45f;
mem_array[39000] = 16'h3e61;
mem_array[39003] = 16'hb256;
mem_array[39002] = 16'h3ef8;
mem_array[39005] = 16'hece2;
mem_array[39004] = 16'h3ef5;
mem_array[39007] = 16'h6504;
mem_array[39006] = 16'h3e6d;
mem_array[39009] = 16'hfac3;
mem_array[39008] = 16'h3ec2;
mem_array[39011] = 16'h40af;
mem_array[39010] = 16'h3e49;
mem_array[39013] = 16'ha6ab;
mem_array[39012] = 16'h3e61;
mem_array[39015] = 16'h61d2;
mem_array[39014] = 16'hbec6;
mem_array[39017] = 16'h3e56;
mem_array[39016] = 16'hbdcd;
mem_array[39019] = 16'hf895;
mem_array[39018] = 16'hbdf3;
mem_array[39021] = 16'hf2ae;
mem_array[39020] = 16'hbcd8;
mem_array[39023] = 16'ha75d;
mem_array[39022] = 16'h3c73;
mem_array[39025] = 16'h3d5a;
mem_array[39024] = 16'hbe1a;
mem_array[39027] = 16'h8bd5;
mem_array[39026] = 16'hbe5d;
mem_array[39029] = 16'h5b07;
mem_array[39028] = 16'h3e97;
mem_array[39031] = 16'hc3f3;
mem_array[39030] = 16'hbd92;
mem_array[39033] = 16'hcfd6;
mem_array[39032] = 16'hbe32;
mem_array[39035] = 16'h2c52;
mem_array[39034] = 16'hbe97;
mem_array[39037] = 16'hc4ce;
mem_array[39036] = 16'hbebc;
mem_array[39039] = 16'h208d;
mem_array[39038] = 16'hbf07;
mem_array[39041] = 16'h4b20;
mem_array[39040] = 16'hbcfb;
mem_array[39043] = 16'hfa2f;
mem_array[39042] = 16'h3c9d;
mem_array[39045] = 16'h4dc8;
mem_array[39044] = 16'hbf39;
mem_array[39047] = 16'h7ce9;
mem_array[39046] = 16'hbd1e;
mem_array[39049] = 16'hf08b;
mem_array[39048] = 16'h3e8f;
mem_array[39051] = 16'h2dd9;
mem_array[39050] = 16'h3f70;
mem_array[39053] = 16'h9273;
mem_array[39052] = 16'h3f03;
mem_array[39055] = 16'h390b;
mem_array[39054] = 16'h3be1;
mem_array[39057] = 16'hdd92;
mem_array[39056] = 16'hbc55;
mem_array[39059] = 16'hc4af;
mem_array[39058] = 16'hbf5f;
mem_array[39061] = 16'h497b;
mem_array[39060] = 16'hbe8d;
mem_array[39063] = 16'hdbf7;
mem_array[39062] = 16'h3ede;
mem_array[39065] = 16'h4277;
mem_array[39064] = 16'h3efc;
mem_array[39067] = 16'h67b9;
mem_array[39066] = 16'h3da7;
mem_array[39069] = 16'h2849;
mem_array[39068] = 16'h3f2b;
mem_array[39071] = 16'ha594;
mem_array[39070] = 16'h3dd8;
mem_array[39073] = 16'h5f72;
mem_array[39072] = 16'h3dd0;
mem_array[39075] = 16'h9722;
mem_array[39074] = 16'h3cc4;
mem_array[39077] = 16'h1f6b;
mem_array[39076] = 16'hbeac;
mem_array[39079] = 16'h924b;
mem_array[39078] = 16'hbf4d;
mem_array[39081] = 16'h658e;
mem_array[39080] = 16'hbbd2;
mem_array[39083] = 16'h8a82;
mem_array[39082] = 16'hbdac;
mem_array[39085] = 16'h20bd;
mem_array[39084] = 16'h3eb6;
mem_array[39087] = 16'hd6ed;
mem_array[39086] = 16'h3d3a;
mem_array[39089] = 16'h3bb9;
mem_array[39088] = 16'h3e81;
mem_array[39091] = 16'had93;
mem_array[39090] = 16'hbdb4;
mem_array[39093] = 16'h1dd8;
mem_array[39092] = 16'hbe39;
mem_array[39095] = 16'he663;
mem_array[39094] = 16'hbc42;
mem_array[39097] = 16'h3d9b;
mem_array[39096] = 16'hbeb2;
mem_array[39099] = 16'h3647;
mem_array[39098] = 16'hbf5d;
mem_array[39101] = 16'hdcb0;
mem_array[39100] = 16'hbec3;
mem_array[39103] = 16'h3ba5;
mem_array[39102] = 16'h3e4c;
mem_array[39105] = 16'h4ff4;
mem_array[39104] = 16'hbfaf;
mem_array[39107] = 16'h1a21;
mem_array[39106] = 16'hbc4a;
mem_array[39109] = 16'h0e28;
mem_array[39108] = 16'h3d4f;
mem_array[39111] = 16'h5a1e;
mem_array[39110] = 16'h3f36;
mem_array[39113] = 16'h72f9;
mem_array[39112] = 16'h3ec9;
mem_array[39115] = 16'hfa2d;
mem_array[39114] = 16'hbbba;
mem_array[39117] = 16'hc933;
mem_array[39116] = 16'hbeab;
mem_array[39119] = 16'hb545;
mem_array[39118] = 16'hbe18;
mem_array[39121] = 16'h0938;
mem_array[39120] = 16'h3e8f;
mem_array[39123] = 16'h2781;
mem_array[39122] = 16'h3ded;
mem_array[39125] = 16'hf71e;
mem_array[39124] = 16'h3e1e;
mem_array[39127] = 16'h9a66;
mem_array[39126] = 16'h3e5f;
mem_array[39129] = 16'h28de;
mem_array[39128] = 16'hbd6c;
mem_array[39131] = 16'hd606;
mem_array[39130] = 16'hbd5e;
mem_array[39133] = 16'h094a;
mem_array[39132] = 16'hba87;
mem_array[39135] = 16'h9ef0;
mem_array[39134] = 16'h3e35;
mem_array[39137] = 16'h6168;
mem_array[39136] = 16'hbb54;
mem_array[39139] = 16'h8602;
mem_array[39138] = 16'hbd6a;
mem_array[39141] = 16'h210d;
mem_array[39140] = 16'hbcf4;
mem_array[39143] = 16'h62b8;
mem_array[39142] = 16'hbd49;
mem_array[39145] = 16'h05f3;
mem_array[39144] = 16'hbd0b;
mem_array[39147] = 16'h1a6f;
mem_array[39146] = 16'hbe87;
mem_array[39149] = 16'h5576;
mem_array[39148] = 16'h3e1c;
mem_array[39151] = 16'h15d0;
mem_array[39150] = 16'h3d44;
mem_array[39153] = 16'hb35a;
mem_array[39152] = 16'h3e2f;
mem_array[39155] = 16'h1e1d;
mem_array[39154] = 16'hbd2b;
mem_array[39157] = 16'hdf9c;
mem_array[39156] = 16'h3d84;
mem_array[39159] = 16'hde49;
mem_array[39158] = 16'hbf23;
mem_array[39161] = 16'h3120;
mem_array[39160] = 16'hbefe;
mem_array[39163] = 16'he592;
mem_array[39162] = 16'h3d8e;
mem_array[39165] = 16'h4ff8;
mem_array[39164] = 16'hbf78;
mem_array[39167] = 16'h73f6;
mem_array[39166] = 16'h3c91;
mem_array[39169] = 16'hc123;
mem_array[39168] = 16'h3cd0;
mem_array[39171] = 16'h05ef;
mem_array[39170] = 16'hbea5;
mem_array[39173] = 16'h916c;
mem_array[39172] = 16'h3dd8;
mem_array[39175] = 16'h1513;
mem_array[39174] = 16'hbe8e;
mem_array[39177] = 16'h67a4;
mem_array[39176] = 16'hbe9f;
mem_array[39179] = 16'hbc94;
mem_array[39178] = 16'hbf17;
mem_array[39181] = 16'hc274;
mem_array[39180] = 16'hbe10;
mem_array[39183] = 16'h6af4;
mem_array[39182] = 16'hbc25;
mem_array[39185] = 16'h96b2;
mem_array[39184] = 16'h3ed2;
mem_array[39187] = 16'h3c3c;
mem_array[39186] = 16'h3e2f;
mem_array[39189] = 16'hccbc;
mem_array[39188] = 16'hbe0b;
mem_array[39191] = 16'hde47;
mem_array[39190] = 16'h3e94;
mem_array[39193] = 16'h24dd;
mem_array[39192] = 16'h3eb4;
mem_array[39195] = 16'hdd0c;
mem_array[39194] = 16'hbdc6;
mem_array[39197] = 16'hdd67;
mem_array[39196] = 16'hbe06;
mem_array[39199] = 16'h23dc;
mem_array[39198] = 16'hbe12;
mem_array[39201] = 16'hdbca;
mem_array[39200] = 16'hbdca;
mem_array[39203] = 16'h9fa2;
mem_array[39202] = 16'hbc19;
mem_array[39205] = 16'hfba6;
mem_array[39204] = 16'hbdee;
mem_array[39207] = 16'hebcc;
mem_array[39206] = 16'hbd8c;
mem_array[39209] = 16'h7d0f;
mem_array[39208] = 16'hbbcc;
mem_array[39211] = 16'hf6fe;
mem_array[39210] = 16'hbdec;
mem_array[39213] = 16'hfec0;
mem_array[39212] = 16'hbdd0;
mem_array[39215] = 16'had40;
mem_array[39214] = 16'hbe58;
mem_array[39217] = 16'h531b;
mem_array[39216] = 16'hbdaa;
mem_array[39219] = 16'h78c6;
mem_array[39218] = 16'hbd83;
mem_array[39221] = 16'hf834;
mem_array[39220] = 16'h3a11;
mem_array[39223] = 16'h2ba0;
mem_array[39222] = 16'hbd59;
mem_array[39225] = 16'h0e5f;
mem_array[39224] = 16'hbe9a;
mem_array[39227] = 16'h5520;
mem_array[39226] = 16'hbe80;
mem_array[39229] = 16'ha32b;
mem_array[39228] = 16'h3deb;
mem_array[39231] = 16'h4eb0;
mem_array[39230] = 16'hbd7e;
mem_array[39233] = 16'h6435;
mem_array[39232] = 16'h3e9b;
mem_array[39235] = 16'he16d;
mem_array[39234] = 16'h3e36;
mem_array[39237] = 16'hf20f;
mem_array[39236] = 16'hbf59;
mem_array[39239] = 16'hd87e;
mem_array[39238] = 16'hbf23;
mem_array[39241] = 16'hff64;
mem_array[39240] = 16'h3c1c;
mem_array[39243] = 16'hd883;
mem_array[39242] = 16'hbdd7;
mem_array[39245] = 16'hed81;
mem_array[39244] = 16'h3e49;
mem_array[39247] = 16'h03d0;
mem_array[39246] = 16'h3ede;
mem_array[39249] = 16'hde12;
mem_array[39248] = 16'hbe53;
mem_array[39251] = 16'hb1f5;
mem_array[39250] = 16'h3e0d;
mem_array[39253] = 16'h87c4;
mem_array[39252] = 16'h3e21;
mem_array[39255] = 16'h8ece;
mem_array[39254] = 16'h3e34;
mem_array[39257] = 16'hd1fa;
mem_array[39256] = 16'hbf04;
mem_array[39259] = 16'h5529;
mem_array[39258] = 16'hbe64;
mem_array[39261] = 16'h78eb;
mem_array[39260] = 16'hbd0b;
mem_array[39263] = 16'hb390;
mem_array[39262] = 16'hbd94;
mem_array[39265] = 16'h470b;
mem_array[39264] = 16'h3e64;
mem_array[39267] = 16'h2728;
mem_array[39266] = 16'hbd3d;
mem_array[39269] = 16'h8278;
mem_array[39268] = 16'hbe2e;
mem_array[39271] = 16'h267f;
mem_array[39270] = 16'hbebe;
mem_array[39273] = 16'h7d13;
mem_array[39272] = 16'hbbd5;
mem_array[39275] = 16'he610;
mem_array[39274] = 16'hbe42;
mem_array[39277] = 16'h790c;
mem_array[39276] = 16'hbc4c;
mem_array[39279] = 16'h7652;
mem_array[39278] = 16'hbda9;
mem_array[39281] = 16'h9e74;
mem_array[39280] = 16'hbca0;
mem_array[39283] = 16'h4fee;
mem_array[39282] = 16'h3cf0;
mem_array[39285] = 16'h769a;
mem_array[39284] = 16'hbf40;
mem_array[39287] = 16'h3442;
mem_array[39286] = 16'hbf0b;
mem_array[39289] = 16'hf478;
mem_array[39288] = 16'hbe23;
mem_array[39291] = 16'h481d;
mem_array[39290] = 16'hbcb8;
mem_array[39293] = 16'heb12;
mem_array[39292] = 16'h3de1;
mem_array[39295] = 16'hf8dd;
mem_array[39294] = 16'h3e90;
mem_array[39297] = 16'h868a;
mem_array[39296] = 16'hbf81;
mem_array[39299] = 16'h3f19;
mem_array[39298] = 16'hbe84;
mem_array[39301] = 16'h3548;
mem_array[39300] = 16'h3e67;
mem_array[39303] = 16'h968f;
mem_array[39302] = 16'hbeb4;
mem_array[39305] = 16'ha6e5;
mem_array[39304] = 16'hbd5f;
mem_array[39307] = 16'he8e0;
mem_array[39306] = 16'h3dcf;
mem_array[39309] = 16'h8aa7;
mem_array[39308] = 16'h3d4a;
mem_array[39311] = 16'ha2d3;
mem_array[39310] = 16'h3d94;
mem_array[39313] = 16'haf46;
mem_array[39312] = 16'h3e04;
mem_array[39315] = 16'h3f72;
mem_array[39314] = 16'hbdac;
mem_array[39317] = 16'h467d;
mem_array[39316] = 16'hbecc;
mem_array[39319] = 16'h1dd3;
mem_array[39318] = 16'hbe02;
mem_array[39321] = 16'h5e13;
mem_array[39320] = 16'hbd27;
mem_array[39323] = 16'h2bc5;
mem_array[39322] = 16'h3c2f;
mem_array[39325] = 16'hb9c6;
mem_array[39324] = 16'hbdd9;
mem_array[39327] = 16'h19c2;
mem_array[39326] = 16'hbe80;
mem_array[39329] = 16'h050c;
mem_array[39328] = 16'h3e02;
mem_array[39331] = 16'h9e06;
mem_array[39330] = 16'hbe5d;
mem_array[39333] = 16'hd9ef;
mem_array[39332] = 16'hbe5c;
mem_array[39335] = 16'h6525;
mem_array[39334] = 16'hbda4;
mem_array[39337] = 16'h6fbc;
mem_array[39336] = 16'hbe20;
mem_array[39339] = 16'hb957;
mem_array[39338] = 16'h3ec5;
mem_array[39341] = 16'h6cac;
mem_array[39340] = 16'hbd0a;
mem_array[39343] = 16'hdc08;
mem_array[39342] = 16'h3e62;
mem_array[39345] = 16'hbcef;
mem_array[39344] = 16'hbf3f;
mem_array[39347] = 16'ha9fb;
mem_array[39346] = 16'hbee3;
mem_array[39349] = 16'h8ea3;
mem_array[39348] = 16'hbd94;
mem_array[39351] = 16'h806d;
mem_array[39350] = 16'hbe08;
mem_array[39353] = 16'h0b7e;
mem_array[39352] = 16'h3e8d;
mem_array[39355] = 16'he30f;
mem_array[39354] = 16'h3e63;
mem_array[39357] = 16'h3dfa;
mem_array[39356] = 16'hbf71;
mem_array[39359] = 16'hf248;
mem_array[39358] = 16'hbe74;
mem_array[39361] = 16'h049d;
mem_array[39360] = 16'hbd34;
mem_array[39363] = 16'hb00a;
mem_array[39362] = 16'h3cfb;
mem_array[39365] = 16'h72b5;
mem_array[39364] = 16'hbcbd;
mem_array[39367] = 16'hf706;
mem_array[39366] = 16'h3c86;
mem_array[39369] = 16'hfc99;
mem_array[39368] = 16'h3e19;
mem_array[39371] = 16'hcd88;
mem_array[39370] = 16'h3d58;
mem_array[39373] = 16'h7dda;
mem_array[39372] = 16'h3d02;
mem_array[39375] = 16'hbf0a;
mem_array[39374] = 16'hbc60;
mem_array[39377] = 16'h0c86;
mem_array[39376] = 16'hbee8;
mem_array[39379] = 16'hffa2;
mem_array[39378] = 16'h3df1;
mem_array[39381] = 16'hb471;
mem_array[39380] = 16'hbc30;
mem_array[39383] = 16'hd604;
mem_array[39382] = 16'h3cbb;
mem_array[39385] = 16'hff11;
mem_array[39384] = 16'hbf0b;
mem_array[39387] = 16'h5baf;
mem_array[39386] = 16'hbee2;
mem_array[39389] = 16'hcdf5;
mem_array[39388] = 16'h3dba;
mem_array[39391] = 16'h8872;
mem_array[39390] = 16'h3d6e;
mem_array[39393] = 16'h55ca;
mem_array[39392] = 16'hbe3f;
mem_array[39395] = 16'hbfc2;
mem_array[39394] = 16'h3d2c;
mem_array[39397] = 16'h5dea;
mem_array[39396] = 16'hbe53;
mem_array[39399] = 16'h0ab5;
mem_array[39398] = 16'h3c74;
mem_array[39401] = 16'h7fdb;
mem_array[39400] = 16'h3c17;
mem_array[39403] = 16'h58f6;
mem_array[39402] = 16'h3cd8;
mem_array[39405] = 16'h22d1;
mem_array[39404] = 16'hbd48;
mem_array[39407] = 16'hd972;
mem_array[39406] = 16'hbdcf;
mem_array[39409] = 16'h4cd1;
mem_array[39408] = 16'hbe29;
mem_array[39411] = 16'h63f8;
mem_array[39410] = 16'hbe82;
mem_array[39413] = 16'hc01d;
mem_array[39412] = 16'h3db1;
mem_array[39415] = 16'h2b62;
mem_array[39414] = 16'h3d15;
mem_array[39417] = 16'hcc7f;
mem_array[39416] = 16'hbefd;
mem_array[39419] = 16'hefa9;
mem_array[39418] = 16'hbee0;
mem_array[39421] = 16'hcf46;
mem_array[39420] = 16'h3eb8;
mem_array[39423] = 16'he246;
mem_array[39422] = 16'h3e61;
mem_array[39425] = 16'h6794;
mem_array[39424] = 16'h3d93;
mem_array[39427] = 16'h807e;
mem_array[39426] = 16'h3d0c;
mem_array[39429] = 16'h62bd;
mem_array[39428] = 16'hbe37;
mem_array[39431] = 16'hcdf1;
mem_array[39430] = 16'hbe4f;
mem_array[39433] = 16'h73c5;
mem_array[39432] = 16'hbd88;
mem_array[39435] = 16'h1c94;
mem_array[39434] = 16'hbdcf;
mem_array[39437] = 16'h3dc2;
mem_array[39436] = 16'hbeab;
mem_array[39439] = 16'h4ac6;
mem_array[39438] = 16'h3d82;
mem_array[39441] = 16'hf357;
mem_array[39440] = 16'hbd4d;
mem_array[39443] = 16'h6cd9;
mem_array[39442] = 16'hbdbe;
mem_array[39445] = 16'ha285;
mem_array[39444] = 16'hbf22;
mem_array[39447] = 16'haab6;
mem_array[39446] = 16'hbed3;
mem_array[39449] = 16'h8401;
mem_array[39448] = 16'hbe2a;
mem_array[39451] = 16'h1780;
mem_array[39450] = 16'h3d8a;
mem_array[39453] = 16'hf654;
mem_array[39452] = 16'hbf08;
mem_array[39455] = 16'h525e;
mem_array[39454] = 16'hbdb5;
mem_array[39457] = 16'h60f4;
mem_array[39456] = 16'hbe25;
mem_array[39459] = 16'h41cd;
mem_array[39458] = 16'hbeeb;
mem_array[39461] = 16'h3c81;
mem_array[39460] = 16'hbe69;
mem_array[39463] = 16'hafe9;
mem_array[39462] = 16'hbdf0;
mem_array[39465] = 16'h1f32;
mem_array[39464] = 16'hbf25;
mem_array[39467] = 16'h9dc8;
mem_array[39466] = 16'hbe1b;
mem_array[39469] = 16'hba38;
mem_array[39468] = 16'hbc38;
mem_array[39471] = 16'h820e;
mem_array[39470] = 16'h3d8a;
mem_array[39473] = 16'h1059;
mem_array[39472] = 16'h3e21;
mem_array[39475] = 16'he139;
mem_array[39474] = 16'hbcf8;
mem_array[39477] = 16'h222b;
mem_array[39476] = 16'hbf59;
mem_array[39479] = 16'hdf7e;
mem_array[39478] = 16'hbedb;
mem_array[39481] = 16'h4208;
mem_array[39480] = 16'h3d3b;
mem_array[39483] = 16'hf6e6;
mem_array[39482] = 16'h3c3c;
mem_array[39485] = 16'h7fae;
mem_array[39484] = 16'h3dd9;
mem_array[39487] = 16'hf64e;
mem_array[39486] = 16'h3e8f;
mem_array[39489] = 16'hc6c8;
mem_array[39488] = 16'hbfce;
mem_array[39491] = 16'hc108;
mem_array[39490] = 16'h3cee;
mem_array[39493] = 16'h50c8;
mem_array[39492] = 16'h3d52;
mem_array[39495] = 16'h3a9d;
mem_array[39494] = 16'hbe64;
mem_array[39497] = 16'h8c1c;
mem_array[39496] = 16'hbdce;
mem_array[39499] = 16'h72af;
mem_array[39498] = 16'hbe3a;
mem_array[39501] = 16'h2d69;
mem_array[39500] = 16'h3d0e;
mem_array[39503] = 16'h3432;
mem_array[39502] = 16'hbcae;
mem_array[39505] = 16'h74ee;
mem_array[39504] = 16'hbeb0;
mem_array[39507] = 16'h3b38;
mem_array[39506] = 16'hbeaa;
mem_array[39509] = 16'h962e;
mem_array[39508] = 16'hbe89;
mem_array[39511] = 16'h029a;
mem_array[39510] = 16'hbe5d;
mem_array[39513] = 16'hb55a;
mem_array[39512] = 16'hbe8f;
mem_array[39515] = 16'h1e35;
mem_array[39514] = 16'h3d95;
mem_array[39517] = 16'h4096;
mem_array[39516] = 16'hbe7d;
mem_array[39519] = 16'hac88;
mem_array[39518] = 16'hbe88;
mem_array[39521] = 16'h4a03;
mem_array[39520] = 16'hbe4f;
mem_array[39523] = 16'hdd32;
mem_array[39522] = 16'hbdff;
mem_array[39525] = 16'h675f;
mem_array[39524] = 16'hbf4b;
mem_array[39527] = 16'h4fd4;
mem_array[39526] = 16'hbd86;
mem_array[39529] = 16'h9735;
mem_array[39528] = 16'hbc72;
mem_array[39531] = 16'h4895;
mem_array[39530] = 16'hbe02;
mem_array[39533] = 16'ha17d;
mem_array[39532] = 16'hbcdb;
mem_array[39535] = 16'h65f5;
mem_array[39534] = 16'h3d05;
mem_array[39537] = 16'h7f39;
mem_array[39536] = 16'hbf94;
mem_array[39539] = 16'haa4b;
mem_array[39538] = 16'hbe99;
mem_array[39541] = 16'h6d91;
mem_array[39540] = 16'hbe1a;
mem_array[39543] = 16'hda74;
mem_array[39542] = 16'h3ea7;
mem_array[39545] = 16'h6ca6;
mem_array[39544] = 16'h3d92;
mem_array[39547] = 16'h7bfa;
mem_array[39546] = 16'hbd91;
mem_array[39549] = 16'h4cfa;
mem_array[39548] = 16'hbf1d;
mem_array[39551] = 16'h4b11;
mem_array[39550] = 16'hbcf7;
mem_array[39553] = 16'hde12;
mem_array[39552] = 16'h3e61;
mem_array[39555] = 16'h19ee;
mem_array[39554] = 16'h3e3a;
mem_array[39557] = 16'h6002;
mem_array[39556] = 16'hbe82;
mem_array[39559] = 16'hc12b;
mem_array[39558] = 16'h3e71;
mem_array[39561] = 16'h5357;
mem_array[39560] = 16'hbdef;
mem_array[39563] = 16'h8872;
mem_array[39562] = 16'hbd0f;
mem_array[39565] = 16'hfedf;
mem_array[39564] = 16'hbf03;
mem_array[39567] = 16'hda2e;
mem_array[39566] = 16'hbead;
mem_array[39569] = 16'h8bc0;
mem_array[39568] = 16'h3e4d;
mem_array[39571] = 16'h4747;
mem_array[39570] = 16'h3e26;
mem_array[39573] = 16'h272b;
mem_array[39572] = 16'hbd47;
mem_array[39575] = 16'h7d41;
mem_array[39574] = 16'hbe6a;
mem_array[39577] = 16'hf773;
mem_array[39576] = 16'hbeeb;
mem_array[39579] = 16'h4c55;
mem_array[39578] = 16'h3e93;
mem_array[39581] = 16'haad3;
mem_array[39580] = 16'hbeb4;
mem_array[39583] = 16'hab6b;
mem_array[39582] = 16'hbe06;
mem_array[39585] = 16'hc338;
mem_array[39584] = 16'hbf1d;
mem_array[39587] = 16'h57fe;
mem_array[39586] = 16'h3b5b;
mem_array[39589] = 16'h2503;
mem_array[39588] = 16'hbe26;
mem_array[39591] = 16'hdd91;
mem_array[39590] = 16'hbc02;
mem_array[39593] = 16'hb4ae;
mem_array[39592] = 16'h3e42;
mem_array[39595] = 16'h6f43;
mem_array[39594] = 16'h3d89;
mem_array[39597] = 16'h3ee2;
mem_array[39596] = 16'hbf1b;
mem_array[39599] = 16'he0dd;
mem_array[39598] = 16'hbdbc;
mem_array[39601] = 16'h5407;
mem_array[39600] = 16'h3ede;
mem_array[39603] = 16'ha475;
mem_array[39602] = 16'h3e82;
mem_array[39605] = 16'h8327;
mem_array[39604] = 16'hbec5;
mem_array[39607] = 16'hef54;
mem_array[39606] = 16'hbdb0;
mem_array[39609] = 16'h91a1;
mem_array[39608] = 16'hbfa9;
mem_array[39611] = 16'hd391;
mem_array[39610] = 16'hbd93;
mem_array[39613] = 16'he29e;
mem_array[39612] = 16'h3d88;
mem_array[39615] = 16'h7090;
mem_array[39614] = 16'hbd7a;
mem_array[39617] = 16'h9238;
mem_array[39616] = 16'hbea2;
mem_array[39619] = 16'h6de3;
mem_array[39618] = 16'h3e5d;
mem_array[39621] = 16'h9ada;
mem_array[39620] = 16'hbd56;
mem_array[39623] = 16'h5e08;
mem_array[39622] = 16'hbde8;
mem_array[39625] = 16'hf73f;
mem_array[39624] = 16'hbfa9;
mem_array[39627] = 16'hff6e;
mem_array[39626] = 16'hbf00;
mem_array[39629] = 16'h3c67;
mem_array[39628] = 16'h3c81;
mem_array[39631] = 16'hcabd;
mem_array[39630] = 16'hbaaa;
mem_array[39633] = 16'h0753;
mem_array[39632] = 16'h3eaa;
mem_array[39635] = 16'hac40;
mem_array[39634] = 16'h3d21;
mem_array[39637] = 16'h4156;
mem_array[39636] = 16'hbed4;
mem_array[39639] = 16'h1b5b;
mem_array[39638] = 16'hbe9f;
mem_array[39641] = 16'h7fd0;
mem_array[39640] = 16'h3ec7;
mem_array[39643] = 16'h72ac;
mem_array[39642] = 16'h3cc6;
mem_array[39645] = 16'h2fba;
mem_array[39644] = 16'hbf04;
mem_array[39647] = 16'h753b;
mem_array[39646] = 16'hbe8a;
mem_array[39649] = 16'he389;
mem_array[39648] = 16'h3e2f;
mem_array[39651] = 16'hb24b;
mem_array[39650] = 16'hbe2a;
mem_array[39653] = 16'h1142;
mem_array[39652] = 16'h3d0e;
mem_array[39655] = 16'h0645;
mem_array[39654] = 16'hbce6;
mem_array[39657] = 16'h98ea;
mem_array[39656] = 16'hbf23;
mem_array[39659] = 16'hd47e;
mem_array[39658] = 16'hbe25;
mem_array[39661] = 16'h76df;
mem_array[39660] = 16'hbeaf;
mem_array[39663] = 16'h8451;
mem_array[39662] = 16'h3eff;
mem_array[39665] = 16'h5c30;
mem_array[39664] = 16'hbeb7;
mem_array[39667] = 16'h7950;
mem_array[39666] = 16'hbb87;
mem_array[39669] = 16'h1063;
mem_array[39668] = 16'hbfe7;
mem_array[39671] = 16'ha8d5;
mem_array[39670] = 16'h3e7a;
mem_array[39673] = 16'h02dc;
mem_array[39672] = 16'hbed4;
mem_array[39675] = 16'haa1a;
mem_array[39674] = 16'hbe9f;
mem_array[39677] = 16'hcbd2;
mem_array[39676] = 16'hbefc;
mem_array[39679] = 16'h239f;
mem_array[39678] = 16'h3e17;
mem_array[39681] = 16'ha567;
mem_array[39680] = 16'hbca9;
mem_array[39683] = 16'h0393;
mem_array[39682] = 16'hbbcc;
mem_array[39685] = 16'he729;
mem_array[39684] = 16'hbf5a;
mem_array[39687] = 16'he140;
mem_array[39686] = 16'hbe0a;
mem_array[39689] = 16'h2fee;
mem_array[39688] = 16'h3eb8;
mem_array[39691] = 16'hebb5;
mem_array[39690] = 16'h3be1;
mem_array[39693] = 16'h9d5c;
mem_array[39692] = 16'h3b8e;
mem_array[39695] = 16'h2a5e;
mem_array[39694] = 16'hbe3f;
mem_array[39697] = 16'h2b03;
mem_array[39696] = 16'hbe88;
mem_array[39699] = 16'h35aa;
mem_array[39698] = 16'hbd67;
mem_array[39701] = 16'haf2b;
mem_array[39700] = 16'h3e7e;
mem_array[39703] = 16'h573a;
mem_array[39702] = 16'hbc9b;
mem_array[39705] = 16'ha028;
mem_array[39704] = 16'hbf3c;
mem_array[39707] = 16'hab8a;
mem_array[39706] = 16'hbcf3;
mem_array[39709] = 16'h0827;
mem_array[39708] = 16'hbe45;
mem_array[39711] = 16'h1e6f;
mem_array[39710] = 16'hbe85;
mem_array[39713] = 16'h017c;
mem_array[39712] = 16'h3da0;
mem_array[39715] = 16'h9e6a;
mem_array[39714] = 16'hbecf;
mem_array[39717] = 16'h2a69;
mem_array[39716] = 16'hbf84;
mem_array[39719] = 16'hc3ca;
mem_array[39718] = 16'hbc4f;
mem_array[39721] = 16'h59d1;
mem_array[39720] = 16'hbec5;
mem_array[39723] = 16'h5b0d;
mem_array[39722] = 16'hbd3c;
mem_array[39725] = 16'hb925;
mem_array[39724] = 16'h3eba;
mem_array[39727] = 16'h49f8;
mem_array[39726] = 16'hbe4c;
mem_array[39729] = 16'hae2e;
mem_array[39728] = 16'hbf0b;
mem_array[39731] = 16'hc6d1;
mem_array[39730] = 16'h3e93;
mem_array[39733] = 16'hb34b;
mem_array[39732] = 16'hbe18;
mem_array[39735] = 16'hece1;
mem_array[39734] = 16'hbef9;
mem_array[39737] = 16'h5cd9;
mem_array[39736] = 16'hbe88;
mem_array[39739] = 16'h7b56;
mem_array[39738] = 16'h3e76;
mem_array[39741] = 16'h9df0;
mem_array[39740] = 16'hbc81;
mem_array[39743] = 16'h4a69;
mem_array[39742] = 16'h3d78;
mem_array[39745] = 16'hc7e5;
mem_array[39744] = 16'hbf4d;
mem_array[39747] = 16'he7b7;
mem_array[39746] = 16'hbeac;
mem_array[39749] = 16'h8bf6;
mem_array[39748] = 16'h3e86;
mem_array[39751] = 16'h8be4;
mem_array[39750] = 16'h3c3a;
mem_array[39753] = 16'h20cc;
mem_array[39752] = 16'h3e0b;
mem_array[39755] = 16'h780b;
mem_array[39754] = 16'h3da5;
mem_array[39757] = 16'h2156;
mem_array[39756] = 16'hbe73;
mem_array[39759] = 16'h50a8;
mem_array[39758] = 16'h3e98;
mem_array[39761] = 16'h8f36;
mem_array[39760] = 16'h3ea7;
mem_array[39763] = 16'h4c2d;
mem_array[39762] = 16'hbf07;
mem_array[39765] = 16'hdaec;
mem_array[39764] = 16'hbec0;
mem_array[39767] = 16'h6dab;
mem_array[39766] = 16'hbe2c;
mem_array[39769] = 16'hf9b7;
mem_array[39768] = 16'hbcb2;
mem_array[39771] = 16'h0a58;
mem_array[39770] = 16'h3dab;
mem_array[39773] = 16'hde60;
mem_array[39772] = 16'hbe2d;
mem_array[39775] = 16'h9f39;
mem_array[39774] = 16'hbc88;
mem_array[39777] = 16'h7abe;
mem_array[39776] = 16'hbe90;
mem_array[39779] = 16'hd030;
mem_array[39778] = 16'h3ed4;
mem_array[39781] = 16'h636e;
mem_array[39780] = 16'h3d8b;
mem_array[39783] = 16'h04e6;
mem_array[39782] = 16'h3bc6;
mem_array[39785] = 16'h5036;
mem_array[39784] = 16'h3e28;
mem_array[39787] = 16'hdb59;
mem_array[39786] = 16'hbf7b;
mem_array[39789] = 16'h3070;
mem_array[39788] = 16'h3db3;
mem_array[39791] = 16'hc40b;
mem_array[39790] = 16'h3bd3;
mem_array[39793] = 16'h2048;
mem_array[39792] = 16'h3e8a;
mem_array[39795] = 16'h1fa9;
mem_array[39794] = 16'hbf3a;
mem_array[39797] = 16'hb4f0;
mem_array[39796] = 16'hbfa4;
mem_array[39799] = 16'h1cfd;
mem_array[39798] = 16'hbee7;
mem_array[39801] = 16'he8f9;
mem_array[39800] = 16'h3ca5;
mem_array[39803] = 16'hc49f;
mem_array[39802] = 16'hbc99;
mem_array[39805] = 16'hc1e9;
mem_array[39804] = 16'hbf5d;
mem_array[39807] = 16'hd504;
mem_array[39806] = 16'hbe5f;
mem_array[39809] = 16'h9062;
mem_array[39808] = 16'h3ed6;
mem_array[39811] = 16'hff54;
mem_array[39810] = 16'h3dc4;
mem_array[39813] = 16'h743c;
mem_array[39812] = 16'h3e82;
mem_array[39815] = 16'h4080;
mem_array[39814] = 16'hbe66;
mem_array[39817] = 16'haccf;
mem_array[39816] = 16'hbe57;
mem_array[39819] = 16'hc8e0;
mem_array[39818] = 16'h3ea1;
mem_array[39821] = 16'h0751;
mem_array[39820] = 16'hbe36;
mem_array[39823] = 16'h4b9c;
mem_array[39822] = 16'hbe86;
mem_array[39825] = 16'h46d5;
mem_array[39824] = 16'hbd16;
mem_array[39827] = 16'hd803;
mem_array[39826] = 16'h3ba1;
mem_array[39829] = 16'h762b;
mem_array[39828] = 16'hbcc2;
mem_array[39831] = 16'h1d10;
mem_array[39830] = 16'hbf8f;
mem_array[39833] = 16'hf667;
mem_array[39832] = 16'hbe03;
mem_array[39835] = 16'h99ee;
mem_array[39834] = 16'h3e6a;
mem_array[39837] = 16'h0b2f;
mem_array[39836] = 16'hbe34;
mem_array[39839] = 16'ha47f;
mem_array[39838] = 16'hbdc8;
mem_array[39841] = 16'h107e;
mem_array[39840] = 16'hbefd;
mem_array[39843] = 16'h76b6;
mem_array[39842] = 16'h3e88;
mem_array[39845] = 16'h253a;
mem_array[39844] = 16'hbe76;
mem_array[39847] = 16'ha29a;
mem_array[39846] = 16'hbf5c;
mem_array[39849] = 16'h743b;
mem_array[39848] = 16'h3eb7;
mem_array[39851] = 16'h97b9;
mem_array[39850] = 16'h3ebd;
mem_array[39853] = 16'h4022;
mem_array[39852] = 16'h3db9;
mem_array[39855] = 16'h9c65;
mem_array[39854] = 16'hbf94;
mem_array[39857] = 16'had36;
mem_array[39856] = 16'hbeea;
mem_array[39859] = 16'h869e;
mem_array[39858] = 16'h3ddf;
mem_array[39861] = 16'h2880;
mem_array[39860] = 16'hb9b0;
mem_array[39863] = 16'h3b34;
mem_array[39862] = 16'hbdcb;
mem_array[39865] = 16'h67a4;
mem_array[39864] = 16'hbf66;
mem_array[39867] = 16'h0080;
mem_array[39866] = 16'h3e04;
mem_array[39869] = 16'ha770;
mem_array[39868] = 16'h3c19;
mem_array[39871] = 16'hf762;
mem_array[39870] = 16'h3e1c;
mem_array[39873] = 16'h0f88;
mem_array[39872] = 16'h3d7a;
mem_array[39875] = 16'hee40;
mem_array[39874] = 16'hbe9b;
mem_array[39877] = 16'h91dc;
mem_array[39876] = 16'hbeb7;
mem_array[39879] = 16'hdeb5;
mem_array[39878] = 16'hbdf2;
mem_array[39881] = 16'h1f6b;
mem_array[39880] = 16'hbed8;
mem_array[39883] = 16'h8380;
mem_array[39882] = 16'h3d26;
mem_array[39885] = 16'h6b28;
mem_array[39884] = 16'hbe9a;
mem_array[39887] = 16'h5837;
mem_array[39886] = 16'hbeca;
mem_array[39889] = 16'hb7ca;
mem_array[39888] = 16'hbccb;
mem_array[39891] = 16'ha41a;
mem_array[39890] = 16'hbf03;
mem_array[39893] = 16'hb770;
mem_array[39892] = 16'h3e8a;
mem_array[39895] = 16'hdbc9;
mem_array[39894] = 16'h3e68;
mem_array[39897] = 16'ha1f3;
mem_array[39896] = 16'hbf68;
mem_array[39899] = 16'h0f44;
mem_array[39898] = 16'h3f15;
mem_array[39901] = 16'hab76;
mem_array[39900] = 16'hbe0d;
mem_array[39903] = 16'hb59d;
mem_array[39902] = 16'hbe05;
mem_array[39905] = 16'h526f;
mem_array[39904] = 16'hbd52;
mem_array[39907] = 16'hd5ec;
mem_array[39906] = 16'hbf58;
mem_array[39909] = 16'h4d20;
mem_array[39908] = 16'h3dec;
mem_array[39911] = 16'h11b4;
mem_array[39910] = 16'hbea5;
mem_array[39913] = 16'h50e9;
mem_array[39912] = 16'h3b79;
mem_array[39915] = 16'h2b30;
mem_array[39914] = 16'hbfc7;
mem_array[39917] = 16'h17a4;
mem_array[39916] = 16'hbe43;
mem_array[39919] = 16'h7341;
mem_array[39918] = 16'hbf01;
mem_array[39921] = 16'he105;
mem_array[39920] = 16'hbd10;
mem_array[39923] = 16'h60c9;
mem_array[39922] = 16'h3d8a;
mem_array[39925] = 16'h4835;
mem_array[39924] = 16'hbf56;
mem_array[39927] = 16'h3bfc;
mem_array[39926] = 16'h3edd;
mem_array[39929] = 16'h5587;
mem_array[39928] = 16'h3e82;
mem_array[39931] = 16'h0900;
mem_array[39930] = 16'h3e28;
mem_array[39933] = 16'h05cf;
mem_array[39932] = 16'h3e3e;
mem_array[39935] = 16'heeab;
mem_array[39934] = 16'h3e9e;
mem_array[39937] = 16'ha523;
mem_array[39936] = 16'hbd81;
mem_array[39939] = 16'hf517;
mem_array[39938] = 16'h3e14;
mem_array[39941] = 16'h696d;
mem_array[39940] = 16'hbe76;
mem_array[39943] = 16'h3896;
mem_array[39942] = 16'hbdd8;
mem_array[39945] = 16'h9344;
mem_array[39944] = 16'hbc84;
mem_array[39947] = 16'h1445;
mem_array[39946] = 16'hbefb;
mem_array[39949] = 16'hac42;
mem_array[39948] = 16'hbe8a;
mem_array[39951] = 16'hedd7;
mem_array[39950] = 16'hbef2;
mem_array[39953] = 16'h65b4;
mem_array[39952] = 16'h3e2f;
mem_array[39955] = 16'h802c;
mem_array[39954] = 16'hbe07;
mem_array[39957] = 16'hca8c;
mem_array[39956] = 16'hbf36;
mem_array[39959] = 16'h2e3c;
mem_array[39958] = 16'h3ee1;
mem_array[39961] = 16'h9fee;
mem_array[39960] = 16'h3d93;
mem_array[39963] = 16'h34d8;
mem_array[39962] = 16'hbeb1;
mem_array[39965] = 16'hf4ab;
mem_array[39964] = 16'h3d5d;
mem_array[39967] = 16'hdf14;
mem_array[39966] = 16'hbef4;
mem_array[39969] = 16'h0b2f;
mem_array[39968] = 16'h3d9b;
mem_array[39971] = 16'h8643;
mem_array[39970] = 16'h3dfc;
mem_array[39973] = 16'h63c6;
mem_array[39972] = 16'hbea8;
mem_array[39975] = 16'h7be3;
mem_array[39974] = 16'hbf8b;
mem_array[39977] = 16'h548a;
mem_array[39976] = 16'hbf88;
mem_array[39979] = 16'h2690;
mem_array[39978] = 16'hbd86;
mem_array[39981] = 16'h9cc4;
mem_array[39980] = 16'hbb00;
mem_array[39983] = 16'hba11;
mem_array[39982] = 16'hbcd5;
mem_array[39985] = 16'h7c3d;
mem_array[39984] = 16'hbf29;
mem_array[39987] = 16'h2ce7;
mem_array[39986] = 16'h3f4f;
mem_array[39989] = 16'h3122;
mem_array[39988] = 16'h3ef3;
mem_array[39991] = 16'h62dc;
mem_array[39990] = 16'h3e7c;
mem_array[39993] = 16'h5243;
mem_array[39992] = 16'h3f2b;
mem_array[39995] = 16'h86c9;
mem_array[39994] = 16'h3db0;
mem_array[39997] = 16'h2351;
mem_array[39996] = 16'hbde1;
mem_array[39999] = 16'hf5ef;
mem_array[39998] = 16'hbf12;
mem_array[40001] = 16'h720c;
mem_array[40000] = 16'h3f4f;
mem_array[40003] = 16'he692;
mem_array[40002] = 16'hbe05;
mem_array[40005] = 16'h6383;
mem_array[40004] = 16'hbf6e;
mem_array[40007] = 16'hb129;
mem_array[40006] = 16'hbebd;
mem_array[40009] = 16'hc194;
mem_array[40008] = 16'h3e62;
mem_array[40011] = 16'h0dfe;
mem_array[40010] = 16'h3e05;
mem_array[40013] = 16'hadde;
mem_array[40012] = 16'h3f45;
mem_array[40015] = 16'h1816;
mem_array[40014] = 16'hbdb0;
mem_array[40017] = 16'h317b;
mem_array[40016] = 16'hbb25;
mem_array[40019] = 16'hef5a;
mem_array[40018] = 16'hbf0f;
mem_array[40021] = 16'hb7d0;
mem_array[40020] = 16'h3dce;
mem_array[40023] = 16'h0896;
mem_array[40022] = 16'hbf90;
mem_array[40025] = 16'h710d;
mem_array[40024] = 16'h3f18;
mem_array[40027] = 16'hfa84;
mem_array[40026] = 16'hbfbf;
mem_array[40029] = 16'hbee7;
mem_array[40028] = 16'hbd6a;
mem_array[40031] = 16'hdf35;
mem_array[40030] = 16'hbe99;
mem_array[40033] = 16'h0616;
mem_array[40032] = 16'hbe02;
mem_array[40035] = 16'h789d;
mem_array[40034] = 16'hbf1b;
mem_array[40037] = 16'hd490;
mem_array[40036] = 16'hbef6;
mem_array[40039] = 16'hcaf6;
mem_array[40038] = 16'hbe03;
mem_array[40041] = 16'h9cc6;
mem_array[40040] = 16'hbd9a;
mem_array[40043] = 16'h7b40;
mem_array[40042] = 16'h3d49;
mem_array[40045] = 16'h1676;
mem_array[40044] = 16'hbf30;
mem_array[40047] = 16'h21ed;
mem_array[40046] = 16'hbe0a;
mem_array[40049] = 16'h182a;
mem_array[40048] = 16'h3f1a;
mem_array[40051] = 16'h27c5;
mem_array[40050] = 16'h3e11;
mem_array[40053] = 16'h9dde;
mem_array[40052] = 16'hbf1d;
mem_array[40055] = 16'h972e;
mem_array[40054] = 16'hbe60;
mem_array[40057] = 16'h5ad5;
mem_array[40056] = 16'hbe42;
mem_array[40059] = 16'h0ee6;
mem_array[40058] = 16'h3d91;
mem_array[40061] = 16'h86d8;
mem_array[40060] = 16'h3f57;
mem_array[40063] = 16'h6a29;
mem_array[40062] = 16'h3e1b;
mem_array[40065] = 16'h119b;
mem_array[40064] = 16'hbf07;
mem_array[40067] = 16'h5426;
mem_array[40066] = 16'h3d8c;
mem_array[40069] = 16'hdebf;
mem_array[40068] = 16'h3cfb;
mem_array[40071] = 16'h00ff;
mem_array[40070] = 16'hbf35;
mem_array[40073] = 16'hfb4d;
mem_array[40072] = 16'h3ece;
mem_array[40075] = 16'hdeb7;
mem_array[40074] = 16'h3d71;
mem_array[40077] = 16'h8dd8;
mem_array[40076] = 16'hbf2a;
mem_array[40079] = 16'hea1f;
mem_array[40078] = 16'hbf20;
mem_array[40081] = 16'h4c4c;
mem_array[40080] = 16'h3f00;
mem_array[40083] = 16'h2549;
mem_array[40082] = 16'hbda8;
mem_array[40085] = 16'h7cdb;
mem_array[40084] = 16'h3f11;
mem_array[40087] = 16'hcabd;
mem_array[40086] = 16'h3e86;
mem_array[40089] = 16'h8bdc;
mem_array[40088] = 16'h3f0a;
mem_array[40091] = 16'h1e82;
mem_array[40090] = 16'hbf90;
mem_array[40093] = 16'hdefe;
mem_array[40092] = 16'hbf28;
mem_array[40095] = 16'hb3f5;
mem_array[40094] = 16'hbea9;
mem_array[40097] = 16'h32c4;
mem_array[40096] = 16'h3d24;
mem_array[40099] = 16'h3d63;
mem_array[40098] = 16'hbe16;
mem_array[40101] = 16'ha703;
mem_array[40100] = 16'hbc2f;
mem_array[40103] = 16'hd8a3;
mem_array[40102] = 16'hbcb0;
mem_array[40105] = 16'h7c3e;
mem_array[40104] = 16'hbee8;
mem_array[40107] = 16'h6b43;
mem_array[40106] = 16'hbec4;
mem_array[40109] = 16'hacc7;
mem_array[40108] = 16'h3f02;
mem_array[40111] = 16'ha3a3;
mem_array[40110] = 16'h3f89;
mem_array[40113] = 16'hef00;
mem_array[40112] = 16'h3fa6;
mem_array[40115] = 16'h6565;
mem_array[40114] = 16'hbeb0;
mem_array[40117] = 16'h9424;
mem_array[40116] = 16'hbf1c;
mem_array[40119] = 16'hf372;
mem_array[40118] = 16'h3c1e;
mem_array[40121] = 16'h3f74;
mem_array[40120] = 16'h3e77;
mem_array[40123] = 16'h9949;
mem_array[40122] = 16'hbb63;
mem_array[40125] = 16'h2c71;
mem_array[40124] = 16'hbe07;
mem_array[40127] = 16'h90b5;
mem_array[40126] = 16'h3f30;
mem_array[40129] = 16'h191c;
mem_array[40128] = 16'hbf1e;
mem_array[40131] = 16'h6e5c;
mem_array[40130] = 16'h3f96;
mem_array[40133] = 16'h7bb2;
mem_array[40132] = 16'h3eb9;
mem_array[40135] = 16'h7a8f;
mem_array[40134] = 16'hbd6e;
mem_array[40137] = 16'h91ef;
mem_array[40136] = 16'hbf3c;
mem_array[40139] = 16'h4cb6;
mem_array[40138] = 16'h3de2;
mem_array[40141] = 16'hd9fa;
mem_array[40140] = 16'h3ea5;
mem_array[40143] = 16'hac55;
mem_array[40142] = 16'hbd9a;
mem_array[40145] = 16'h0051;
mem_array[40144] = 16'h3d16;
mem_array[40147] = 16'h9d8a;
mem_array[40146] = 16'h3f24;
mem_array[40149] = 16'hc9ca;
mem_array[40148] = 16'h3ddd;
mem_array[40151] = 16'h82b0;
mem_array[40150] = 16'hbef6;
mem_array[40153] = 16'h198c;
mem_array[40152] = 16'hbf26;
mem_array[40155] = 16'hda1e;
mem_array[40154] = 16'hbe76;
mem_array[40157] = 16'h3501;
mem_array[40156] = 16'hbe28;
mem_array[40159] = 16'hfe70;
mem_array[40158] = 16'h3dd6;
mem_array[40161] = 16'hb70b;
mem_array[40160] = 16'h3bff;
mem_array[40163] = 16'h5849;
mem_array[40162] = 16'h3a32;
mem_array[40165] = 16'h90c1;
mem_array[40164] = 16'h3f1c;
mem_array[40167] = 16'h5b40;
mem_array[40166] = 16'hbfb2;
mem_array[40169] = 16'haaa0;
mem_array[40168] = 16'h3d2a;
mem_array[40171] = 16'hb821;
mem_array[40170] = 16'h3f97;
mem_array[40173] = 16'h02f9;
mem_array[40172] = 16'h3f67;
mem_array[40175] = 16'h8011;
mem_array[40174] = 16'h3f4e;
mem_array[40177] = 16'h09b0;
mem_array[40176] = 16'h3ea6;
mem_array[40179] = 16'hc49e;
mem_array[40178] = 16'h3ec9;
mem_array[40181] = 16'h14e4;
mem_array[40180] = 16'h3f7d;
mem_array[40183] = 16'h5993;
mem_array[40182] = 16'hbf1c;
mem_array[40185] = 16'h4d14;
mem_array[40184] = 16'hbda2;
mem_array[40187] = 16'h7a6d;
mem_array[40186] = 16'h3f8b;
mem_array[40189] = 16'h5151;
mem_array[40188] = 16'hbf10;
mem_array[40191] = 16'ha5b4;
mem_array[40190] = 16'h3f04;
mem_array[40193] = 16'h7634;
mem_array[40192] = 16'hbe10;
mem_array[40195] = 16'h6692;
mem_array[40194] = 16'h3eb0;
mem_array[40197] = 16'h2b91;
mem_array[40196] = 16'hbef0;
mem_array[40199] = 16'h43d6;
mem_array[40198] = 16'h3eea;
mem_array[40201] = 16'h9734;
mem_array[40200] = 16'h3f8a;
mem_array[40203] = 16'h052c;
mem_array[40202] = 16'h3d1a;
mem_array[40205] = 16'h27d3;
mem_array[40204] = 16'hbea5;
mem_array[40207] = 16'h75cd;
mem_array[40206] = 16'h3efc;
mem_array[40209] = 16'h50ad;
mem_array[40208] = 16'h3e2b;
mem_array[40211] = 16'ha1f3;
mem_array[40210] = 16'h3e8d;
mem_array[40213] = 16'h115c;
mem_array[40212] = 16'hbe11;
mem_array[40215] = 16'ha63c;
mem_array[40214] = 16'hbe58;
mem_array[40217] = 16'hd76f;
mem_array[40216] = 16'hbe9e;
mem_array[40219] = 16'h1525;
mem_array[40218] = 16'h3f8a;
mem_array[40221] = 16'h40d9;
mem_array[40220] = 16'hbd34;
mem_array[40223] = 16'hbe60;
mem_array[40222] = 16'h3d52;
mem_array[40225] = 16'h6812;
mem_array[40224] = 16'h3f71;
mem_array[40227] = 16'h0704;
mem_array[40226] = 16'hbfc1;
mem_array[40229] = 16'ha7e3;
mem_array[40228] = 16'hbe6c;
mem_array[40231] = 16'hae87;
mem_array[40230] = 16'h3e4b;
mem_array[40233] = 16'h9423;
mem_array[40232] = 16'h3ed9;
mem_array[40235] = 16'hfba4;
mem_array[40234] = 16'h3f59;
mem_array[40237] = 16'h6fbd;
mem_array[40236] = 16'hbeac;
mem_array[40239] = 16'h8d9f;
mem_array[40238] = 16'h3f44;
mem_array[40241] = 16'h3b2d;
mem_array[40240] = 16'h3f1d;
mem_array[40243] = 16'h11ce;
mem_array[40242] = 16'hbf24;
mem_array[40245] = 16'h7047;
mem_array[40244] = 16'hbcd4;
mem_array[40247] = 16'h255c;
mem_array[40246] = 16'h3d50;
mem_array[40249] = 16'h673a;
mem_array[40248] = 16'hbd49;
mem_array[40251] = 16'he722;
mem_array[40250] = 16'hbc5d;
mem_array[40253] = 16'he51b;
mem_array[40252] = 16'hbf31;
mem_array[40255] = 16'h41a1;
mem_array[40254] = 16'h3ce1;
mem_array[40257] = 16'h8e4c;
mem_array[40256] = 16'hbf30;
mem_array[40259] = 16'h7f30;
mem_array[40258] = 16'h3f58;
mem_array[40261] = 16'h7d2e;
mem_array[40260] = 16'hba9f;
mem_array[40263] = 16'h1ac4;
mem_array[40262] = 16'h3d29;
mem_array[40265] = 16'hc2b7;
mem_array[40264] = 16'hbc95;
mem_array[40267] = 16'hc442;
mem_array[40266] = 16'hbd8a;
mem_array[40269] = 16'h39e1;
mem_array[40268] = 16'h3d27;
mem_array[40271] = 16'h1a35;
mem_array[40270] = 16'hbdb4;
mem_array[40273] = 16'h617e;
mem_array[40272] = 16'hbd45;
mem_array[40275] = 16'hc70a;
mem_array[40274] = 16'h3d4f;
mem_array[40277] = 16'hee90;
mem_array[40276] = 16'hbd3f;
mem_array[40279] = 16'h68eb;
mem_array[40278] = 16'hbddd;
mem_array[40281] = 16'h296d;
mem_array[40280] = 16'h3d80;
mem_array[40283] = 16'hc93f;
mem_array[40282] = 16'h3dd0;
mem_array[40285] = 16'ha80d;
mem_array[40284] = 16'h3d18;
mem_array[40287] = 16'hfe8e;
mem_array[40286] = 16'h3d8f;
mem_array[40289] = 16'h4792;
mem_array[40288] = 16'h3cc4;
mem_array[40291] = 16'heaaf;
mem_array[40290] = 16'hbce4;
mem_array[40293] = 16'h6388;
mem_array[40292] = 16'h3d50;
mem_array[40295] = 16'hb4db;
mem_array[40294] = 16'h3daa;
mem_array[40297] = 16'h00d4;
mem_array[40296] = 16'hbbdd;
mem_array[40299] = 16'h948e;
mem_array[40298] = 16'h3dbc;
mem_array[40301] = 16'h5dd4;
mem_array[40300] = 16'h3c81;
mem_array[40303] = 16'h7199;
mem_array[40302] = 16'h3a38;
mem_array[40305] = 16'he2cd;
mem_array[40304] = 16'hbcee;
mem_array[40307] = 16'h0fbe;
mem_array[40306] = 16'h3d83;
mem_array[40309] = 16'heb11;
mem_array[40308] = 16'h3d09;
mem_array[40311] = 16'hc6c5;
mem_array[40310] = 16'h3c68;
mem_array[40313] = 16'h7c1e;
mem_array[40312] = 16'hbd84;
mem_array[40315] = 16'h80a1;
mem_array[40314] = 16'hbbe2;
mem_array[40317] = 16'hdb18;
mem_array[40316] = 16'h3dad;
mem_array[40319] = 16'hff72;
mem_array[40318] = 16'h3d8e;
mem_array[40321] = 16'he43b;
mem_array[40320] = 16'h3d0c;
mem_array[40323] = 16'ha17b;
mem_array[40322] = 16'h3d38;
mem_array[40325] = 16'h8fd5;
mem_array[40324] = 16'hbd80;
mem_array[40327] = 16'haa69;
mem_array[40326] = 16'h3c84;
mem_array[40329] = 16'hb832;
mem_array[40328] = 16'hbd89;
mem_array[40331] = 16'h452b;
mem_array[40330] = 16'hbcd3;
mem_array[40333] = 16'h342e;
mem_array[40332] = 16'h3dda;
mem_array[40335] = 16'hee17;
mem_array[40334] = 16'hbd39;
mem_array[40337] = 16'ha90d;
mem_array[40336] = 16'hbc8e;
mem_array[40339] = 16'he3d9;
mem_array[40338] = 16'h3c51;
mem_array[40341] = 16'ha0b9;
mem_array[40340] = 16'hbd63;
mem_array[40343] = 16'hc4ba;
mem_array[40342] = 16'h3d81;
mem_array[40345] = 16'h79af;
mem_array[40344] = 16'hb997;
mem_array[40347] = 16'h30c4;
mem_array[40346] = 16'h3d56;
mem_array[40349] = 16'h5ac3;
mem_array[40348] = 16'hbb96;
mem_array[40351] = 16'h91f6;
mem_array[40350] = 16'hbc9f;
mem_array[40353] = 16'h1b7e;
mem_array[40352] = 16'hbd75;
mem_array[40355] = 16'hcf28;
mem_array[40354] = 16'hbdc4;
mem_array[40357] = 16'hef1f;
mem_array[40356] = 16'h3d95;
mem_array[40359] = 16'h6333;
mem_array[40358] = 16'hbdae;
mem_array[40361] = 16'hc166;
mem_array[40360] = 16'h3b1e;
mem_array[40363] = 16'h9c1a;
mem_array[40362] = 16'hbd30;
mem_array[40365] = 16'h8f2f;
mem_array[40364] = 16'hbcb4;
mem_array[40367] = 16'h0e84;
mem_array[40366] = 16'hbc88;
mem_array[40369] = 16'h4af1;
mem_array[40368] = 16'hbc53;
mem_array[40371] = 16'hbca0;
mem_array[40370] = 16'hbdb5;
mem_array[40373] = 16'hc968;
mem_array[40372] = 16'h3b8d;
mem_array[40375] = 16'h8a16;
mem_array[40374] = 16'hbb8b;
mem_array[40377] = 16'h29b5;
mem_array[40376] = 16'hbd20;
mem_array[40379] = 16'h50e7;
mem_array[40378] = 16'h3daa;
mem_array[40381] = 16'h6c75;
mem_array[40380] = 16'h3cc3;
mem_array[40383] = 16'hdcdf;
mem_array[40382] = 16'hbd1b;
mem_array[40385] = 16'h1cb2;
mem_array[40384] = 16'hbcbd;
mem_array[40387] = 16'h1a3e;
mem_array[40386] = 16'hbc9a;
mem_array[40389] = 16'h59db;
mem_array[40388] = 16'h3cc5;
mem_array[40391] = 16'h8ac2;
mem_array[40390] = 16'hbb64;
mem_array[40393] = 16'h5ff5;
mem_array[40392] = 16'h3ca5;
mem_array[40395] = 16'h830e;
mem_array[40394] = 16'h3c59;
mem_array[40397] = 16'h9208;
mem_array[40396] = 16'h3d9b;
mem_array[40399] = 16'h2204;
mem_array[40398] = 16'h3d32;
mem_array[40401] = 16'hffe2;
mem_array[40400] = 16'hbb5b;
mem_array[40403] = 16'h99eb;
mem_array[40402] = 16'h3bbb;
mem_array[40405] = 16'h8b17;
mem_array[40404] = 16'h3daa;
mem_array[40407] = 16'h6299;
mem_array[40406] = 16'h3cf7;
mem_array[40409] = 16'hdd2f;
mem_array[40408] = 16'h3de6;
mem_array[40411] = 16'ha977;
mem_array[40410] = 16'h3d1e;
mem_array[40413] = 16'h2898;
mem_array[40412] = 16'h3d4f;
mem_array[40415] = 16'h3f99;
mem_array[40414] = 16'hbc8c;
mem_array[40417] = 16'ha969;
mem_array[40416] = 16'h3dbf;
mem_array[40419] = 16'h2a98;
mem_array[40418] = 16'h3db3;
mem_array[40421] = 16'hbae1;
mem_array[40420] = 16'hbccf;
mem_array[40423] = 16'h60c3;
mem_array[40422] = 16'hbc0a;
mem_array[40425] = 16'h665e;
mem_array[40424] = 16'h3dd9;
mem_array[40427] = 16'h0530;
mem_array[40426] = 16'hbdc2;
mem_array[40429] = 16'h2a2a;
mem_array[40428] = 16'hba5b;
mem_array[40431] = 16'h799e;
mem_array[40430] = 16'h3d68;
mem_array[40433] = 16'h8580;
mem_array[40432] = 16'h3dde;
mem_array[40435] = 16'h6e21;
mem_array[40434] = 16'hbd26;
mem_array[40437] = 16'hff11;
mem_array[40436] = 16'hbd08;
mem_array[40439] = 16'h5d3a;
mem_array[40438] = 16'hbd77;
mem_array[40441] = 16'h7ac8;
mem_array[40440] = 16'hbc16;
mem_array[40443] = 16'h3fc3;
mem_array[40442] = 16'h3da1;
mem_array[40445] = 16'ha35b;
mem_array[40444] = 16'h3ec6;
mem_array[40447] = 16'he8fa;
mem_array[40446] = 16'h3c0d;
mem_array[40449] = 16'hdbbe;
mem_array[40448] = 16'h3e46;
mem_array[40451] = 16'hf30d;
mem_array[40450] = 16'hbe9c;
mem_array[40453] = 16'h96e3;
mem_array[40452] = 16'h3eb5;
mem_array[40455] = 16'h80c7;
mem_array[40454] = 16'h3db1;
mem_array[40457] = 16'h28c7;
mem_array[40456] = 16'h3c69;
mem_array[40459] = 16'h2fc2;
mem_array[40458] = 16'h3cb1;
mem_array[40461] = 16'he1f4;
mem_array[40460] = 16'hbce7;
mem_array[40463] = 16'h4369;
mem_array[40462] = 16'h3d46;
mem_array[40465] = 16'h1e70;
mem_array[40464] = 16'h3d58;
mem_array[40467] = 16'h9893;
mem_array[40466] = 16'h3e3a;
mem_array[40469] = 16'h2863;
mem_array[40468] = 16'hbe0e;
mem_array[40471] = 16'h06bc;
mem_array[40470] = 16'hbe01;
mem_array[40473] = 16'he5b8;
mem_array[40472] = 16'hbd6d;
mem_array[40475] = 16'h3a17;
mem_array[40474] = 16'h3d35;
mem_array[40477] = 16'hf984;
mem_array[40476] = 16'hbdad;
mem_array[40479] = 16'h6a04;
mem_array[40478] = 16'hbd7d;
mem_array[40481] = 16'h77c2;
mem_array[40480] = 16'hbdf1;
mem_array[40483] = 16'h3af2;
mem_array[40482] = 16'hbe5e;
mem_array[40485] = 16'h1fb1;
mem_array[40484] = 16'hbd4c;
mem_array[40487] = 16'hd146;
mem_array[40486] = 16'hbe90;
mem_array[40489] = 16'h1e9a;
mem_array[40488] = 16'hbd3c;
mem_array[40491] = 16'h9884;
mem_array[40490] = 16'hbdfd;
mem_array[40493] = 16'h8f77;
mem_array[40492] = 16'h3e54;
mem_array[40495] = 16'hf513;
mem_array[40494] = 16'hbc90;
mem_array[40497] = 16'h6c64;
mem_array[40496] = 16'hbe3c;
mem_array[40499] = 16'ha69a;
mem_array[40498] = 16'hbe76;
mem_array[40501] = 16'h4b73;
mem_array[40500] = 16'hbef9;
mem_array[40503] = 16'h6839;
mem_array[40502] = 16'hbe0e;
mem_array[40505] = 16'hfb95;
mem_array[40504] = 16'hbeb0;
mem_array[40507] = 16'hceba;
mem_array[40506] = 16'h3dcd;
mem_array[40509] = 16'h464d;
mem_array[40508] = 16'hbec1;
mem_array[40511] = 16'h14d7;
mem_array[40510] = 16'hbe31;
mem_array[40513] = 16'h79b2;
mem_array[40512] = 16'h3e94;
mem_array[40515] = 16'h37ed;
mem_array[40514] = 16'hbeb1;
mem_array[40517] = 16'h740d;
mem_array[40516] = 16'hbf24;
mem_array[40519] = 16'h42d7;
mem_array[40518] = 16'hbc50;
mem_array[40521] = 16'h5056;
mem_array[40520] = 16'hbc0f;
mem_array[40523] = 16'h23f2;
mem_array[40522] = 16'hbca1;
mem_array[40525] = 16'heaa8;
mem_array[40524] = 16'hbea5;
mem_array[40527] = 16'hdf47;
mem_array[40526] = 16'hbfab;
mem_array[40529] = 16'h8eee;
mem_array[40528] = 16'hbdae;
mem_array[40531] = 16'hae26;
mem_array[40530] = 16'hbf89;
mem_array[40533] = 16'h5317;
mem_array[40532] = 16'hbe89;
mem_array[40535] = 16'h3301;
mem_array[40534] = 16'h3cbf;
mem_array[40537] = 16'hcd74;
mem_array[40536] = 16'hbf2e;
mem_array[40539] = 16'h8ad0;
mem_array[40538] = 16'hbcae;
mem_array[40541] = 16'hc2d9;
mem_array[40540] = 16'hbe48;
mem_array[40543] = 16'h89ab;
mem_array[40542] = 16'h3ea1;
mem_array[40545] = 16'hde23;
mem_array[40544] = 16'hbe43;
mem_array[40547] = 16'h18cd;
mem_array[40546] = 16'hbeda;
mem_array[40549] = 16'h7234;
mem_array[40548] = 16'h3f25;
mem_array[40551] = 16'he043;
mem_array[40550] = 16'h3d3c;
mem_array[40553] = 16'h90f7;
mem_array[40552] = 16'h3f7c;
mem_array[40555] = 16'h03bd;
mem_array[40554] = 16'h3c21;
mem_array[40557] = 16'hadaa;
mem_array[40556] = 16'h3e6c;
mem_array[40559] = 16'h7c7f;
mem_array[40558] = 16'hbcdf;
mem_array[40561] = 16'hacb4;
mem_array[40560] = 16'hbe19;
mem_array[40563] = 16'h8047;
mem_array[40562] = 16'hbea5;
mem_array[40565] = 16'h9a21;
mem_array[40564] = 16'hbed2;
mem_array[40567] = 16'hf54e;
mem_array[40566] = 16'h3ef7;
mem_array[40569] = 16'h8697;
mem_array[40568] = 16'h3eed;
mem_array[40571] = 16'h8d3a;
mem_array[40570] = 16'h3f76;
mem_array[40573] = 16'haf98;
mem_array[40572] = 16'h3db9;
mem_array[40575] = 16'ha5e0;
mem_array[40574] = 16'hbde7;
mem_array[40577] = 16'h5678;
mem_array[40576] = 16'hbf46;
mem_array[40579] = 16'he5f4;
mem_array[40578] = 16'h3d3d;
mem_array[40581] = 16'h37f7;
mem_array[40580] = 16'hbb22;
mem_array[40583] = 16'hccaa;
mem_array[40582] = 16'h3d7f;
mem_array[40585] = 16'ha38e;
mem_array[40584] = 16'hbf70;
mem_array[40587] = 16'h0f95;
mem_array[40586] = 16'hbf8d;
mem_array[40589] = 16'head6;
mem_array[40588] = 16'h3e36;
mem_array[40591] = 16'hcb57;
mem_array[40590] = 16'hbedf;
mem_array[40593] = 16'hac7e;
mem_array[40592] = 16'hbf0b;
mem_array[40595] = 16'h4efe;
mem_array[40594] = 16'hbec4;
mem_array[40597] = 16'h78ef;
mem_array[40596] = 16'hc002;
mem_array[40599] = 16'hf0c4;
mem_array[40598] = 16'hbea0;
mem_array[40601] = 16'hd67d;
mem_array[40600] = 16'hbef4;
mem_array[40603] = 16'h1548;
mem_array[40602] = 16'h3f1a;
mem_array[40605] = 16'h0b9e;
mem_array[40604] = 16'hbcc6;
mem_array[40607] = 16'h58ba;
mem_array[40606] = 16'hbf10;
mem_array[40609] = 16'h4444;
mem_array[40608] = 16'h3f55;
mem_array[40611] = 16'hd0fb;
mem_array[40610] = 16'h3f5a;
mem_array[40613] = 16'h375a;
mem_array[40612] = 16'h3ed2;
mem_array[40615] = 16'hf92c;
mem_array[40614] = 16'hbe3f;
mem_array[40617] = 16'hfd6c;
mem_array[40616] = 16'hbd07;
mem_array[40619] = 16'ha2ca;
mem_array[40618] = 16'h3d56;
mem_array[40621] = 16'h7b6b;
mem_array[40620] = 16'h3eca;
mem_array[40623] = 16'h9657;
mem_array[40622] = 16'h3e81;
mem_array[40625] = 16'h7df5;
mem_array[40624] = 16'hbea4;
mem_array[40627] = 16'h699c;
mem_array[40626] = 16'h3f68;
mem_array[40629] = 16'hbd58;
mem_array[40628] = 16'h3eb7;
mem_array[40631] = 16'h3a3a;
mem_array[40630] = 16'h3f4f;
mem_array[40633] = 16'heb4a;
mem_array[40632] = 16'hbdca;
mem_array[40635] = 16'hdf2f;
mem_array[40634] = 16'h3da0;
mem_array[40637] = 16'h44ea;
mem_array[40636] = 16'hbf93;
mem_array[40639] = 16'h94a2;
mem_array[40638] = 16'hbe99;
mem_array[40641] = 16'hbeed;
mem_array[40640] = 16'h3dbc;
mem_array[40643] = 16'h843f;
mem_array[40642] = 16'hbdd1;
mem_array[40645] = 16'ha671;
mem_array[40644] = 16'hbf70;
mem_array[40647] = 16'h9b7f;
mem_array[40646] = 16'hbf78;
mem_array[40649] = 16'ha07a;
mem_array[40648] = 16'h3e84;
mem_array[40651] = 16'ha3a0;
mem_array[40650] = 16'hbd03;
mem_array[40653] = 16'h04bb;
mem_array[40652] = 16'hbee2;
mem_array[40655] = 16'h4373;
mem_array[40654] = 16'h3e4a;
mem_array[40657] = 16'hae47;
mem_array[40656] = 16'hbf15;
mem_array[40659] = 16'hed45;
mem_array[40658] = 16'h3db7;
mem_array[40661] = 16'hcddd;
mem_array[40660] = 16'hbec5;
mem_array[40663] = 16'h444e;
mem_array[40662] = 16'h3f1a;
mem_array[40665] = 16'he0b4;
mem_array[40664] = 16'hbd2b;
mem_array[40667] = 16'h6628;
mem_array[40666] = 16'hbf05;
mem_array[40669] = 16'h6cfe;
mem_array[40668] = 16'h3ec6;
mem_array[40671] = 16'h1849;
mem_array[40670] = 16'h3f69;
mem_array[40673] = 16'h8e59;
mem_array[40672] = 16'h3ec4;
mem_array[40675] = 16'h7c00;
mem_array[40674] = 16'h3ed9;
mem_array[40677] = 16'h6bc7;
mem_array[40676] = 16'hbf34;
mem_array[40679] = 16'hd781;
mem_array[40678] = 16'h3f02;
mem_array[40681] = 16'hc3b3;
mem_array[40680] = 16'hbd3b;
mem_array[40683] = 16'hbe78;
mem_array[40682] = 16'h3e01;
mem_array[40685] = 16'h8cc4;
mem_array[40684] = 16'hbe93;
mem_array[40687] = 16'h3f45;
mem_array[40686] = 16'h3ef1;
mem_array[40689] = 16'hd16e;
mem_array[40688] = 16'h3f0b;
mem_array[40691] = 16'ha2ce;
mem_array[40690] = 16'h3d12;
mem_array[40693] = 16'hecdb;
mem_array[40692] = 16'h3e43;
mem_array[40695] = 16'h0886;
mem_array[40694] = 16'hbe87;
mem_array[40697] = 16'h71e2;
mem_array[40696] = 16'hbf1c;
mem_array[40699] = 16'ha1c7;
mem_array[40698] = 16'h3f55;
mem_array[40701] = 16'h2541;
mem_array[40700] = 16'hbc3a;
mem_array[40703] = 16'h3539;
mem_array[40702] = 16'h3d92;
mem_array[40705] = 16'he7ee;
mem_array[40704] = 16'hbfaf;
mem_array[40707] = 16'h7bf8;
mem_array[40706] = 16'hbfc8;
mem_array[40709] = 16'h564d;
mem_array[40708] = 16'hbe2a;
mem_array[40711] = 16'h8fb7;
mem_array[40710] = 16'hbc0c;
mem_array[40713] = 16'h72b7;
mem_array[40712] = 16'hbf44;
mem_array[40715] = 16'hce22;
mem_array[40714] = 16'h3f3a;
mem_array[40717] = 16'hf847;
mem_array[40716] = 16'hbf77;
mem_array[40719] = 16'h7d20;
mem_array[40718] = 16'hbd3b;
mem_array[40721] = 16'h7747;
mem_array[40720] = 16'h3dcf;
mem_array[40723] = 16'h2e19;
mem_array[40722] = 16'h3eeb;
mem_array[40725] = 16'hbdb5;
mem_array[40724] = 16'h3dbe;
mem_array[40727] = 16'h8e59;
mem_array[40726] = 16'h3ea4;
mem_array[40729] = 16'h33e6;
mem_array[40728] = 16'h3eab;
mem_array[40731] = 16'h293b;
mem_array[40730] = 16'hbd59;
mem_array[40733] = 16'hbf6d;
mem_array[40732] = 16'h3ce1;
mem_array[40735] = 16'h6833;
mem_array[40734] = 16'hbdc0;
mem_array[40737] = 16'hb942;
mem_array[40736] = 16'hbf57;
mem_array[40739] = 16'h4119;
mem_array[40738] = 16'hbf36;
mem_array[40741] = 16'h1e6d;
mem_array[40740] = 16'hbf02;
mem_array[40743] = 16'h2bbb;
mem_array[40742] = 16'h3ed2;
mem_array[40745] = 16'he199;
mem_array[40744] = 16'hbe58;
mem_array[40747] = 16'h7924;
mem_array[40746] = 16'h3da5;
mem_array[40749] = 16'heeaf;
mem_array[40748] = 16'h3f17;
mem_array[40751] = 16'hbf44;
mem_array[40750] = 16'hbdce;
mem_array[40753] = 16'h2907;
mem_array[40752] = 16'h3d22;
mem_array[40755] = 16'hd756;
mem_array[40754] = 16'h3d77;
mem_array[40757] = 16'h827b;
mem_array[40756] = 16'hbefb;
mem_array[40759] = 16'h552c;
mem_array[40758] = 16'hbf12;
mem_array[40761] = 16'h2be8;
mem_array[40760] = 16'h3d3c;
mem_array[40763] = 16'hb80f;
mem_array[40762] = 16'hbc1f;
mem_array[40765] = 16'h967f;
mem_array[40764] = 16'hbfa6;
mem_array[40767] = 16'hf886;
mem_array[40766] = 16'hbf54;
mem_array[40769] = 16'h7b26;
mem_array[40768] = 16'hbe10;
mem_array[40771] = 16'h1d49;
mem_array[40770] = 16'hbe60;
mem_array[40773] = 16'h4cf6;
mem_array[40772] = 16'hbf3f;
mem_array[40775] = 16'h1e17;
mem_array[40774] = 16'h3ed2;
mem_array[40777] = 16'h997e;
mem_array[40776] = 16'h3de3;
mem_array[40779] = 16'hff95;
mem_array[40778] = 16'hbf6f;
mem_array[40781] = 16'h1339;
mem_array[40780] = 16'hbee4;
mem_array[40783] = 16'h6628;
mem_array[40782] = 16'h3eef;
mem_array[40785] = 16'hccc0;
mem_array[40784] = 16'h3db2;
mem_array[40787] = 16'h1fd9;
mem_array[40786] = 16'hbe24;
mem_array[40789] = 16'hc351;
mem_array[40788] = 16'h3e55;
mem_array[40791] = 16'heaab;
mem_array[40790] = 16'hbe22;
mem_array[40793] = 16'h6fd5;
mem_array[40792] = 16'h3de5;
mem_array[40795] = 16'h2d3e;
mem_array[40794] = 16'hbe8d;
mem_array[40797] = 16'h426c;
mem_array[40796] = 16'hbf48;
mem_array[40799] = 16'h6a48;
mem_array[40798] = 16'hbf0c;
mem_array[40801] = 16'h5bf5;
mem_array[40800] = 16'hbee7;
mem_array[40803] = 16'hbe2e;
mem_array[40802] = 16'h3e37;
mem_array[40805] = 16'hd0c9;
mem_array[40804] = 16'h3e4b;
mem_array[40807] = 16'h12ce;
mem_array[40806] = 16'h3b3b;
mem_array[40809] = 16'hda5b;
mem_array[40808] = 16'h3f13;
mem_array[40811] = 16'h45ac;
mem_array[40810] = 16'hbe65;
mem_array[40813] = 16'hd859;
mem_array[40812] = 16'h3e7b;
mem_array[40815] = 16'h87bf;
mem_array[40814] = 16'h3e8e;
mem_array[40817] = 16'hb0a5;
mem_array[40816] = 16'hbec6;
mem_array[40819] = 16'h9bdb;
mem_array[40818] = 16'hbf99;
mem_array[40821] = 16'hf370;
mem_array[40820] = 16'h3bbc;
mem_array[40823] = 16'ha85e;
mem_array[40822] = 16'h3c14;
mem_array[40825] = 16'h3439;
mem_array[40824] = 16'hbf76;
mem_array[40827] = 16'hd838;
mem_array[40826] = 16'hbf88;
mem_array[40829] = 16'ha831;
mem_array[40828] = 16'hbf2f;
mem_array[40831] = 16'h45db;
mem_array[40830] = 16'hbdd6;
mem_array[40833] = 16'h6338;
mem_array[40832] = 16'hbf21;
mem_array[40835] = 16'hdee7;
mem_array[40834] = 16'hbe89;
mem_array[40837] = 16'h1915;
mem_array[40836] = 16'hbd05;
mem_array[40839] = 16'hb518;
mem_array[40838] = 16'hbe53;
mem_array[40841] = 16'h85be;
mem_array[40840] = 16'hbeeb;
mem_array[40843] = 16'hf8a6;
mem_array[40842] = 16'h3e00;
mem_array[40845] = 16'hd5c9;
mem_array[40844] = 16'hbe08;
mem_array[40847] = 16'h6787;
mem_array[40846] = 16'hbd6e;
mem_array[40849] = 16'ha79c;
mem_array[40848] = 16'h3e26;
mem_array[40851] = 16'hf804;
mem_array[40850] = 16'h3ebf;
mem_array[40853] = 16'hbcd0;
mem_array[40852] = 16'h3e03;
mem_array[40855] = 16'h891a;
mem_array[40854] = 16'hbebe;
mem_array[40857] = 16'ha5c2;
mem_array[40856] = 16'hbf0a;
mem_array[40859] = 16'h025b;
mem_array[40858] = 16'hbe05;
mem_array[40861] = 16'h3a80;
mem_array[40860] = 16'hbbca;
mem_array[40863] = 16'h86e2;
mem_array[40862] = 16'hbe95;
mem_array[40865] = 16'h9a8d;
mem_array[40864] = 16'h3e3e;
mem_array[40867] = 16'h34bb;
mem_array[40866] = 16'h3b4d;
mem_array[40869] = 16'h0efe;
mem_array[40868] = 16'hbcfd;
mem_array[40871] = 16'hd68d;
mem_array[40870] = 16'h3ea6;
mem_array[40873] = 16'h80bd;
mem_array[40872] = 16'h3def;
mem_array[40875] = 16'hcc63;
mem_array[40874] = 16'hbf43;
mem_array[40877] = 16'h9fd2;
mem_array[40876] = 16'hbf7a;
mem_array[40879] = 16'h07db;
mem_array[40878] = 16'hbe0e;
mem_array[40881] = 16'h9bd6;
mem_array[40880] = 16'h3dbf;
mem_array[40883] = 16'h0b92;
mem_array[40882] = 16'hbd77;
mem_array[40885] = 16'h2f63;
mem_array[40884] = 16'hbf7e;
mem_array[40887] = 16'hfc15;
mem_array[40886] = 16'hbf56;
mem_array[40889] = 16'h7f96;
mem_array[40888] = 16'hbf08;
mem_array[40891] = 16'h6ab8;
mem_array[40890] = 16'hbeea;
mem_array[40893] = 16'h5c95;
mem_array[40892] = 16'h3ebc;
mem_array[40895] = 16'he703;
mem_array[40894] = 16'h3ec4;
mem_array[40897] = 16'hcf70;
mem_array[40896] = 16'hbec5;
mem_array[40899] = 16'h8bc9;
mem_array[40898] = 16'h3ea7;
mem_array[40901] = 16'hdcf0;
mem_array[40900] = 16'hbda4;
mem_array[40903] = 16'h8fb9;
mem_array[40902] = 16'h3cd9;
mem_array[40905] = 16'h32c3;
mem_array[40904] = 16'hbfa0;
mem_array[40907] = 16'he2bb;
mem_array[40906] = 16'hbe81;
mem_array[40909] = 16'h74f7;
mem_array[40908] = 16'hbd19;
mem_array[40911] = 16'hd4de;
mem_array[40910] = 16'h3d97;
mem_array[40913] = 16'h17aa;
mem_array[40912] = 16'h3e4d;
mem_array[40915] = 16'hcfac;
mem_array[40914] = 16'h3e2a;
mem_array[40917] = 16'he677;
mem_array[40916] = 16'hbf1a;
mem_array[40919] = 16'heb4d;
mem_array[40918] = 16'hbed4;
mem_array[40921] = 16'h3a72;
mem_array[40920] = 16'hbdb1;
mem_array[40923] = 16'h8b37;
mem_array[40922] = 16'h3de5;
mem_array[40925] = 16'h12f8;
mem_array[40924] = 16'hbecf;
mem_array[40927] = 16'h4bbc;
mem_array[40926] = 16'h3e00;
mem_array[40929] = 16'hbc42;
mem_array[40928] = 16'h3dcb;
mem_array[40931] = 16'h03d3;
mem_array[40930] = 16'h3d30;
mem_array[40933] = 16'h9534;
mem_array[40932] = 16'h3efe;
mem_array[40935] = 16'ha29a;
mem_array[40934] = 16'hbf1c;
mem_array[40937] = 16'hc83b;
mem_array[40936] = 16'hbf61;
mem_array[40939] = 16'habed;
mem_array[40938] = 16'hbe71;
mem_array[40941] = 16'h070b;
mem_array[40940] = 16'hbd00;
mem_array[40943] = 16'h054e;
mem_array[40942] = 16'h3c14;
mem_array[40945] = 16'hdef2;
mem_array[40944] = 16'hbf7f;
mem_array[40947] = 16'ha7dd;
mem_array[40946] = 16'hbef4;
mem_array[40949] = 16'h5d97;
mem_array[40948] = 16'hbf05;
mem_array[40951] = 16'hc641;
mem_array[40950] = 16'hbcda;
mem_array[40953] = 16'h311b;
mem_array[40952] = 16'hbe93;
mem_array[40955] = 16'h3423;
mem_array[40954] = 16'hbe02;
mem_array[40957] = 16'h6726;
mem_array[40956] = 16'hbdec;
mem_array[40959] = 16'h02d8;
mem_array[40958] = 16'h3d25;
mem_array[40961] = 16'h99b7;
mem_array[40960] = 16'hbe2a;
mem_array[40963] = 16'hda7d;
mem_array[40962] = 16'h3dd3;
mem_array[40965] = 16'hd4e7;
mem_array[40964] = 16'hbf98;
mem_array[40967] = 16'hec50;
mem_array[40966] = 16'h3e06;
mem_array[40969] = 16'h7e33;
mem_array[40968] = 16'h3cf2;
mem_array[40971] = 16'h11a9;
mem_array[40970] = 16'hbcad;
mem_array[40973] = 16'h8a6c;
mem_array[40972] = 16'h3d4e;
mem_array[40975] = 16'h6697;
mem_array[40974] = 16'h3c00;
mem_array[40977] = 16'h4458;
mem_array[40976] = 16'hbf35;
mem_array[40979] = 16'h6fae;
mem_array[40978] = 16'hbd5c;
mem_array[40981] = 16'h97d3;
mem_array[40980] = 16'hbde2;
mem_array[40983] = 16'h248b;
mem_array[40982] = 16'h3e5b;
mem_array[40985] = 16'h3cec;
mem_array[40984] = 16'hbd4e;
mem_array[40987] = 16'h4523;
mem_array[40986] = 16'hbe6b;
mem_array[40989] = 16'h7a3b;
mem_array[40988] = 16'h3eef;
mem_array[40991] = 16'h5726;
mem_array[40990] = 16'hbe61;
mem_array[40993] = 16'hdba3;
mem_array[40992] = 16'h3e82;
mem_array[40995] = 16'h822a;
mem_array[40994] = 16'hbf1f;
mem_array[40997] = 16'hf08e;
mem_array[40996] = 16'hbed8;
mem_array[40999] = 16'hf43b;
mem_array[40998] = 16'hbe55;
mem_array[41001] = 16'h54ae;
mem_array[41000] = 16'h3c08;
mem_array[41003] = 16'h52ce;
mem_array[41002] = 16'h3d57;
mem_array[41005] = 16'h3bd2;
mem_array[41004] = 16'hbf42;
mem_array[41007] = 16'h31d7;
mem_array[41006] = 16'hbee9;
mem_array[41009] = 16'h4ad3;
mem_array[41008] = 16'hbd65;
mem_array[41011] = 16'h2152;
mem_array[41010] = 16'hbd3a;
mem_array[41013] = 16'hdffd;
mem_array[41012] = 16'hbd2b;
mem_array[41015] = 16'h7f4a;
mem_array[41014] = 16'hbe43;
mem_array[41017] = 16'h6bfc;
mem_array[41016] = 16'hbe11;
mem_array[41019] = 16'h3758;
mem_array[41018] = 16'h3ebd;
mem_array[41021] = 16'hfa16;
mem_array[41020] = 16'hbc8e;
mem_array[41023] = 16'heb07;
mem_array[41022] = 16'hbd86;
mem_array[41025] = 16'h4df1;
mem_array[41024] = 16'hbfc1;
mem_array[41027] = 16'h9c10;
mem_array[41026] = 16'hbc8b;
mem_array[41029] = 16'h5632;
mem_array[41028] = 16'h3e40;
mem_array[41031] = 16'h9608;
mem_array[41030] = 16'h3f06;
mem_array[41033] = 16'h2bff;
mem_array[41032] = 16'h3e1b;
mem_array[41035] = 16'h68ae;
mem_array[41034] = 16'h3e7f;
mem_array[41037] = 16'h3c5c;
mem_array[41036] = 16'hbe02;
mem_array[41039] = 16'h4d83;
mem_array[41038] = 16'hbd4a;
mem_array[41041] = 16'haea4;
mem_array[41040] = 16'h3edd;
mem_array[41043] = 16'h76d8;
mem_array[41042] = 16'hbba5;
mem_array[41045] = 16'h36ec;
mem_array[41044] = 16'h3e0f;
mem_array[41047] = 16'h5bd3;
mem_array[41046] = 16'h3ead;
mem_array[41049] = 16'h6237;
mem_array[41048] = 16'h3f38;
mem_array[41051] = 16'h9fee;
mem_array[41050] = 16'hbd1c;
mem_array[41053] = 16'hebae;
mem_array[41052] = 16'hbe83;
mem_array[41055] = 16'h77de;
mem_array[41054] = 16'hbf32;
mem_array[41057] = 16'h1f0e;
mem_array[41056] = 16'hbdef;
mem_array[41059] = 16'h6b84;
mem_array[41058] = 16'hbe92;
mem_array[41061] = 16'h2000;
mem_array[41060] = 16'hbd3b;
mem_array[41063] = 16'h30cd;
mem_array[41062] = 16'h3c00;
mem_array[41065] = 16'he9a7;
mem_array[41064] = 16'hbe90;
mem_array[41067] = 16'h575a;
mem_array[41066] = 16'hbf43;
mem_array[41069] = 16'h6ef9;
mem_array[41068] = 16'h3d3d;
mem_array[41071] = 16'ha9f2;
mem_array[41070] = 16'hbe44;
mem_array[41073] = 16'h84d0;
mem_array[41072] = 16'h3e92;
mem_array[41075] = 16'h2fbb;
mem_array[41074] = 16'h3e01;
mem_array[41077] = 16'h3691;
mem_array[41076] = 16'hbe8e;
mem_array[41079] = 16'h1221;
mem_array[41078] = 16'h3dd8;
mem_array[41081] = 16'he0b4;
mem_array[41080] = 16'hbd6e;
mem_array[41083] = 16'h7177;
mem_array[41082] = 16'hbe5f;
mem_array[41085] = 16'h10f2;
mem_array[41084] = 16'hbfbf;
mem_array[41087] = 16'he19d;
mem_array[41086] = 16'h3da6;
mem_array[41089] = 16'h0f80;
mem_array[41088] = 16'hbe89;
mem_array[41091] = 16'h7576;
mem_array[41090] = 16'h3e59;
mem_array[41093] = 16'he356;
mem_array[41092] = 16'h3e59;
mem_array[41095] = 16'h63e1;
mem_array[41094] = 16'h3de1;
mem_array[41097] = 16'h0e56;
mem_array[41096] = 16'h3e0d;
mem_array[41099] = 16'hebdb;
mem_array[41098] = 16'hbede;
mem_array[41101] = 16'ha592;
mem_array[41100] = 16'h3e0e;
mem_array[41103] = 16'h9e87;
mem_array[41102] = 16'hbc8c;
mem_array[41105] = 16'h6d22;
mem_array[41104] = 16'hbe5d;
mem_array[41107] = 16'h2225;
mem_array[41106] = 16'h3df4;
mem_array[41109] = 16'h6522;
mem_array[41108] = 16'hbec8;
mem_array[41111] = 16'h5518;
mem_array[41110] = 16'hbe47;
mem_array[41113] = 16'h35bd;
mem_array[41112] = 16'h3e9a;
mem_array[41115] = 16'h68d6;
mem_array[41114] = 16'hbf26;
mem_array[41117] = 16'hae22;
mem_array[41116] = 16'hbf23;
mem_array[41119] = 16'h93e3;
mem_array[41118] = 16'hbf4c;
mem_array[41121] = 16'h7019;
mem_array[41120] = 16'h3ce2;
mem_array[41123] = 16'h2b40;
mem_array[41122] = 16'hbdcf;
mem_array[41125] = 16'h4e60;
mem_array[41124] = 16'hbe3c;
mem_array[41127] = 16'h7d5b;
mem_array[41126] = 16'hbf3f;
mem_array[41129] = 16'h6a40;
mem_array[41128] = 16'h3d24;
mem_array[41131] = 16'haa4b;
mem_array[41130] = 16'hbe24;
mem_array[41133] = 16'h8715;
mem_array[41132] = 16'h3e0e;
mem_array[41135] = 16'hd46d;
mem_array[41134] = 16'h3eb2;
mem_array[41137] = 16'he3cf;
mem_array[41136] = 16'hbeb7;
mem_array[41139] = 16'h243a;
mem_array[41138] = 16'h3e2e;
mem_array[41141] = 16'hfc9a;
mem_array[41140] = 16'hbbe1;
mem_array[41143] = 16'h9a58;
mem_array[41142] = 16'h3dd0;
mem_array[41145] = 16'h3e44;
mem_array[41144] = 16'hbf71;
mem_array[41147] = 16'hba35;
mem_array[41146] = 16'hbcc9;
mem_array[41149] = 16'h2fbe;
mem_array[41148] = 16'h3dcf;
mem_array[41151] = 16'h64dc;
mem_array[41150] = 16'hbd52;
mem_array[41153] = 16'h63ab;
mem_array[41152] = 16'h3e90;
mem_array[41155] = 16'h278e;
mem_array[41154] = 16'h3e24;
mem_array[41157] = 16'h2afa;
mem_array[41156] = 16'hbed4;
mem_array[41159] = 16'h57ea;
mem_array[41158] = 16'h3e9b;
mem_array[41161] = 16'h2f8c;
mem_array[41160] = 16'h3eae;
mem_array[41163] = 16'h8f5e;
mem_array[41162] = 16'h3e47;
mem_array[41165] = 16'hc4f2;
mem_array[41164] = 16'h3e67;
mem_array[41167] = 16'hd976;
mem_array[41166] = 16'h3cc8;
mem_array[41169] = 16'h982c;
mem_array[41168] = 16'hbf8b;
mem_array[41171] = 16'h2107;
mem_array[41170] = 16'hbe0a;
mem_array[41173] = 16'h19f6;
mem_array[41172] = 16'h3e6d;
mem_array[41175] = 16'hc801;
mem_array[41174] = 16'hbef7;
mem_array[41177] = 16'h1ef5;
mem_array[41176] = 16'hbecc;
mem_array[41179] = 16'h3770;
mem_array[41178] = 16'hbf41;
mem_array[41181] = 16'h535d;
mem_array[41180] = 16'hbcc1;
mem_array[41183] = 16'hdd07;
mem_array[41182] = 16'h3d73;
mem_array[41185] = 16'h6028;
mem_array[41184] = 16'hbf3b;
mem_array[41187] = 16'hd941;
mem_array[41186] = 16'hbf3b;
mem_array[41189] = 16'haffd;
mem_array[41188] = 16'hbe91;
mem_array[41191] = 16'he793;
mem_array[41190] = 16'hbd3a;
mem_array[41193] = 16'hc406;
mem_array[41192] = 16'h3de2;
mem_array[41195] = 16'h6007;
mem_array[41194] = 16'h3ead;
mem_array[41197] = 16'hdc0a;
mem_array[41196] = 16'hbf01;
mem_array[41199] = 16'haf34;
mem_array[41198] = 16'h3e2c;
mem_array[41201] = 16'hdf26;
mem_array[41200] = 16'hbcfc;
mem_array[41203] = 16'h8005;
mem_array[41202] = 16'h3e22;
mem_array[41205] = 16'h4f30;
mem_array[41204] = 16'hbfe9;
mem_array[41207] = 16'hc942;
mem_array[41206] = 16'h3d8c;
mem_array[41209] = 16'hb21c;
mem_array[41208] = 16'hbdde;
mem_array[41211] = 16'hb083;
mem_array[41210] = 16'hbd42;
mem_array[41213] = 16'h8014;
mem_array[41212] = 16'h3e90;
mem_array[41215] = 16'h080c;
mem_array[41214] = 16'h3e2c;
mem_array[41217] = 16'h9e61;
mem_array[41216] = 16'hbf73;
mem_array[41219] = 16'hc2fb;
mem_array[41218] = 16'h3da7;
mem_array[41221] = 16'h2fc7;
mem_array[41220] = 16'h3fb1;
mem_array[41223] = 16'h174d;
mem_array[41222] = 16'hbe37;
mem_array[41225] = 16'h96e6;
mem_array[41224] = 16'h3e3d;
mem_array[41227] = 16'h908c;
mem_array[41226] = 16'h3d01;
mem_array[41229] = 16'h0a08;
mem_array[41228] = 16'hbfd4;
mem_array[41231] = 16'h95c4;
mem_array[41230] = 16'h3c72;
mem_array[41233] = 16'h4e8d;
mem_array[41232] = 16'h3e3f;
mem_array[41235] = 16'hde82;
mem_array[41234] = 16'hbebc;
mem_array[41237] = 16'hcd47;
mem_array[41236] = 16'hbc71;
mem_array[41239] = 16'ha5cf;
mem_array[41238] = 16'hbe93;
mem_array[41241] = 16'hd86d;
mem_array[41240] = 16'hbd8c;
mem_array[41243] = 16'h9783;
mem_array[41242] = 16'hbd6c;
mem_array[41245] = 16'hc194;
mem_array[41244] = 16'hbf9b;
mem_array[41247] = 16'h73ba;
mem_array[41246] = 16'hbf3a;
mem_array[41249] = 16'h56ec;
mem_array[41248] = 16'hbc92;
mem_array[41251] = 16'hcff0;
mem_array[41250] = 16'hbc62;
mem_array[41253] = 16'h6be6;
mem_array[41252] = 16'h3d83;
mem_array[41255] = 16'h0e87;
mem_array[41254] = 16'hbea5;
mem_array[41257] = 16'h6a43;
mem_array[41256] = 16'hbe8a;
mem_array[41259] = 16'hdf77;
mem_array[41258] = 16'h3d9b;
mem_array[41261] = 16'hcedd;
mem_array[41260] = 16'hbec4;
mem_array[41263] = 16'h1fb9;
mem_array[41262] = 16'h3d87;
mem_array[41265] = 16'h48f9;
mem_array[41264] = 16'hbfb4;
mem_array[41267] = 16'h783c;
mem_array[41266] = 16'hbc42;
mem_array[41269] = 16'h424e;
mem_array[41268] = 16'hbd6a;
mem_array[41271] = 16'h08fc;
mem_array[41270] = 16'hbde9;
mem_array[41273] = 16'hc77c;
mem_array[41272] = 16'h3de6;
mem_array[41275] = 16'h64ff;
mem_array[41274] = 16'h3c8c;
mem_array[41277] = 16'h456e;
mem_array[41276] = 16'hbefd;
mem_array[41279] = 16'hf416;
mem_array[41278] = 16'hbe8c;
mem_array[41281] = 16'h5d2e;
mem_array[41280] = 16'hbe62;
mem_array[41283] = 16'hea67;
mem_array[41282] = 16'h3e0d;
mem_array[41285] = 16'habff;
mem_array[41284] = 16'hbdc9;
mem_array[41287] = 16'hd4a1;
mem_array[41286] = 16'hbe5f;
mem_array[41289] = 16'hf6c8;
mem_array[41288] = 16'hbfcd;
mem_array[41291] = 16'h94f6;
mem_array[41290] = 16'hbf05;
mem_array[41293] = 16'had4e;
mem_array[41292] = 16'h3ca0;
mem_array[41295] = 16'hce88;
mem_array[41294] = 16'hbf67;
mem_array[41297] = 16'ha67e;
mem_array[41296] = 16'h3e1b;
mem_array[41299] = 16'h9b97;
mem_array[41298] = 16'h3e01;
mem_array[41301] = 16'hc168;
mem_array[41300] = 16'h3cd2;
mem_array[41303] = 16'h3e63;
mem_array[41302] = 16'hbc7a;
mem_array[41305] = 16'h06de;
mem_array[41304] = 16'hbfff;
mem_array[41307] = 16'h1d5f;
mem_array[41306] = 16'hbf34;
mem_array[41309] = 16'h0111;
mem_array[41308] = 16'hbf11;
mem_array[41311] = 16'hafe1;
mem_array[41310] = 16'hbcd5;
mem_array[41313] = 16'h4570;
mem_array[41312] = 16'h3e4d;
mem_array[41315] = 16'h51e4;
mem_array[41314] = 16'h3ee2;
mem_array[41317] = 16'h9a46;
mem_array[41316] = 16'hbe5d;
mem_array[41319] = 16'he944;
mem_array[41318] = 16'h3e1a;
mem_array[41321] = 16'haf88;
mem_array[41320] = 16'hbdaf;
mem_array[41323] = 16'hb40d;
mem_array[41322] = 16'hbe30;
mem_array[41325] = 16'ha7d2;
mem_array[41324] = 16'hbdc7;
mem_array[41327] = 16'h8eb4;
mem_array[41326] = 16'h3e3d;
mem_array[41329] = 16'hbbde;
mem_array[41328] = 16'hbe15;
mem_array[41331] = 16'h2c03;
mem_array[41330] = 16'hbecf;
mem_array[41333] = 16'h74d6;
mem_array[41332] = 16'h3e1b;
mem_array[41335] = 16'h3180;
mem_array[41334] = 16'hbe98;
mem_array[41337] = 16'hc955;
mem_array[41336] = 16'hbf14;
mem_array[41339] = 16'haa1c;
mem_array[41338] = 16'hbdc0;
mem_array[41341] = 16'h15c6;
mem_array[41340] = 16'hbf8e;
mem_array[41343] = 16'h6c69;
mem_array[41342] = 16'h3e7c;
mem_array[41345] = 16'hb56c;
mem_array[41344] = 16'hbed1;
mem_array[41347] = 16'habcb;
mem_array[41346] = 16'hbed7;
mem_array[41349] = 16'h6b35;
mem_array[41348] = 16'hbfb0;
mem_array[41351] = 16'hf559;
mem_array[41350] = 16'hbe6d;
mem_array[41353] = 16'hb3b8;
mem_array[41352] = 16'hbd91;
mem_array[41355] = 16'h9a81;
mem_array[41354] = 16'hbe2d;
mem_array[41357] = 16'ha115;
mem_array[41356] = 16'h3eb4;
mem_array[41359] = 16'hc464;
mem_array[41358] = 16'h3e71;
mem_array[41361] = 16'hd157;
mem_array[41360] = 16'hbc56;
mem_array[41363] = 16'h0477;
mem_array[41362] = 16'h3d2f;
mem_array[41365] = 16'hc84e;
mem_array[41364] = 16'hbff2;
mem_array[41367] = 16'hec33;
mem_array[41366] = 16'hbe71;
mem_array[41369] = 16'hd431;
mem_array[41368] = 16'hbd6a;
mem_array[41371] = 16'h6828;
mem_array[41370] = 16'hbe9e;
mem_array[41373] = 16'h3359;
mem_array[41372] = 16'h3e07;
mem_array[41375] = 16'h43aa;
mem_array[41374] = 16'h3e12;
mem_array[41377] = 16'h4b94;
mem_array[41376] = 16'hbe03;
mem_array[41379] = 16'ha3ca;
mem_array[41378] = 16'hbdf0;
mem_array[41381] = 16'h10ca;
mem_array[41380] = 16'hbec4;
mem_array[41383] = 16'h4dea;
mem_array[41382] = 16'h3d68;
mem_array[41385] = 16'h7e4a;
mem_array[41384] = 16'hbfe2;
mem_array[41387] = 16'h9912;
mem_array[41386] = 16'h3daf;
mem_array[41389] = 16'hf448;
mem_array[41388] = 16'h3e87;
mem_array[41391] = 16'hfd60;
mem_array[41390] = 16'hbecb;
mem_array[41393] = 16'h4804;
mem_array[41392] = 16'h3e91;
mem_array[41395] = 16'hd2b3;
mem_array[41394] = 16'hbd8d;
mem_array[41397] = 16'hb97f;
mem_array[41396] = 16'hbee6;
mem_array[41399] = 16'h4955;
mem_array[41398] = 16'hbf08;
mem_array[41401] = 16'h27d3;
mem_array[41400] = 16'hbfb3;
mem_array[41403] = 16'h8ea3;
mem_array[41402] = 16'hbe8b;
mem_array[41405] = 16'h5c16;
mem_array[41404] = 16'hbaae;
mem_array[41407] = 16'h7b1c;
mem_array[41406] = 16'hbf80;
mem_array[41409] = 16'h85c8;
mem_array[41408] = 16'hbfd1;
mem_array[41411] = 16'h7813;
mem_array[41410] = 16'hbe72;
mem_array[41413] = 16'he172;
mem_array[41412] = 16'hbe9d;
mem_array[41415] = 16'h8926;
mem_array[41414] = 16'hbe70;
mem_array[41417] = 16'hbeca;
mem_array[41416] = 16'h3dd6;
mem_array[41419] = 16'h58de;
mem_array[41418] = 16'hbf19;
mem_array[41421] = 16'h5848;
mem_array[41420] = 16'hbd8e;
mem_array[41423] = 16'hff0f;
mem_array[41422] = 16'h3d2d;
mem_array[41425] = 16'hcfda;
mem_array[41424] = 16'hc00e;
mem_array[41427] = 16'hd5ea;
mem_array[41426] = 16'hbee5;
mem_array[41429] = 16'hacc0;
mem_array[41428] = 16'hbe26;
mem_array[41431] = 16'hd1f5;
mem_array[41430] = 16'h38d5;
mem_array[41433] = 16'hef31;
mem_array[41432] = 16'h3ed0;
mem_array[41435] = 16'h3322;
mem_array[41434] = 16'h3e9f;
mem_array[41437] = 16'h14a6;
mem_array[41436] = 16'hbdff;
mem_array[41439] = 16'hf187;
mem_array[41438] = 16'hbf1e;
mem_array[41441] = 16'ha0ab;
mem_array[41440] = 16'h3cbe;
mem_array[41443] = 16'hc899;
mem_array[41442] = 16'h3e89;
mem_array[41445] = 16'hc723;
mem_array[41444] = 16'hbfa3;
mem_array[41447] = 16'h4d3c;
mem_array[41446] = 16'h3d2f;
mem_array[41449] = 16'h02c6;
mem_array[41448] = 16'hbf2f;
mem_array[41451] = 16'h25c3;
mem_array[41450] = 16'hbf43;
mem_array[41453] = 16'h932c;
mem_array[41452] = 16'h3e4b;
mem_array[41455] = 16'h31d4;
mem_array[41454] = 16'h3e06;
mem_array[41457] = 16'h0ded;
mem_array[41456] = 16'hbeb2;
mem_array[41459] = 16'hedbf;
mem_array[41458] = 16'h3f0c;
mem_array[41461] = 16'h7641;
mem_array[41460] = 16'hbfac;
mem_array[41463] = 16'h7fd2;
mem_array[41462] = 16'hbe03;
mem_array[41465] = 16'hcbae;
mem_array[41464] = 16'hbe4d;
mem_array[41467] = 16'h40e3;
mem_array[41466] = 16'hbfa6;
mem_array[41469] = 16'h3e5c;
mem_array[41468] = 16'hbf81;
mem_array[41471] = 16'hcd8a;
mem_array[41470] = 16'hbe00;
mem_array[41473] = 16'ha659;
mem_array[41472] = 16'hbe3d;
mem_array[41475] = 16'h7bbe;
mem_array[41474] = 16'hbf9b;
mem_array[41477] = 16'hf8ad;
mem_array[41476] = 16'hbf44;
mem_array[41479] = 16'hf4de;
mem_array[41478] = 16'hbf17;
mem_array[41481] = 16'haf94;
mem_array[41480] = 16'h3d70;
mem_array[41483] = 16'h70c9;
mem_array[41482] = 16'hbd16;
mem_array[41485] = 16'h56d0;
mem_array[41484] = 16'hbff3;
mem_array[41487] = 16'hf13e;
mem_array[41486] = 16'hbf1c;
mem_array[41489] = 16'hb9d6;
mem_array[41488] = 16'h3f05;
mem_array[41491] = 16'h9e8e;
mem_array[41490] = 16'h3e28;
mem_array[41493] = 16'hdd37;
mem_array[41492] = 16'h3e5e;
mem_array[41495] = 16'h597a;
mem_array[41494] = 16'hbe72;
mem_array[41497] = 16'h7852;
mem_array[41496] = 16'hbc85;
mem_array[41499] = 16'h93c5;
mem_array[41498] = 16'hbee4;
mem_array[41501] = 16'hede5;
mem_array[41500] = 16'hbd80;
mem_array[41503] = 16'h9ebd;
mem_array[41502] = 16'h3e84;
mem_array[41505] = 16'hb234;
mem_array[41504] = 16'hbf92;
mem_array[41507] = 16'h200b;
mem_array[41506] = 16'h3be4;
mem_array[41509] = 16'heb18;
mem_array[41508] = 16'hbf18;
mem_array[41511] = 16'hbd18;
mem_array[41510] = 16'hbf5f;
mem_array[41513] = 16'h1707;
mem_array[41512] = 16'h3da8;
mem_array[41515] = 16'hd55e;
mem_array[41514] = 16'h3dcf;
mem_array[41517] = 16'h203c;
mem_array[41516] = 16'hbec2;
mem_array[41519] = 16'h1ec9;
mem_array[41518] = 16'h3eb1;
mem_array[41521] = 16'h32e5;
mem_array[41520] = 16'hbf85;
mem_array[41523] = 16'hcb40;
mem_array[41522] = 16'h3e7b;
mem_array[41525] = 16'h1d07;
mem_array[41524] = 16'hbe33;
mem_array[41527] = 16'heabe;
mem_array[41526] = 16'hbfbc;
mem_array[41529] = 16'h06a9;
mem_array[41528] = 16'hbe67;
mem_array[41531] = 16'hc212;
mem_array[41530] = 16'hbf77;
mem_array[41533] = 16'ha43b;
mem_array[41532] = 16'hbda4;
mem_array[41535] = 16'he32f;
mem_array[41534] = 16'hbf60;
mem_array[41537] = 16'hbe69;
mem_array[41536] = 16'hbe9b;
mem_array[41539] = 16'h750d;
mem_array[41538] = 16'hbf2b;
mem_array[41541] = 16'h3626;
mem_array[41540] = 16'hbc76;
mem_array[41543] = 16'h982e;
mem_array[41542] = 16'hbc48;
mem_array[41545] = 16'hd23a;
mem_array[41544] = 16'hc000;
mem_array[41547] = 16'h0ede;
mem_array[41546] = 16'hbebb;
mem_array[41549] = 16'hf2ba;
mem_array[41548] = 16'h3e53;
mem_array[41551] = 16'hb865;
mem_array[41550] = 16'hbc22;
mem_array[41553] = 16'h989d;
mem_array[41552] = 16'h3e8f;
mem_array[41555] = 16'hbd28;
mem_array[41554] = 16'h3daf;
mem_array[41557] = 16'ha151;
mem_array[41556] = 16'h3e45;
mem_array[41559] = 16'h1aaa;
mem_array[41558] = 16'hbde2;
mem_array[41561] = 16'hfb0d;
mem_array[41560] = 16'h3e4a;
mem_array[41563] = 16'h681f;
mem_array[41562] = 16'h3e04;
mem_array[41565] = 16'h7a7a;
mem_array[41564] = 16'hbf40;
mem_array[41567] = 16'h5171;
mem_array[41566] = 16'hbeca;
mem_array[41569] = 16'h7f57;
mem_array[41568] = 16'h3e54;
mem_array[41571] = 16'h72ce;
mem_array[41570] = 16'hbdcd;
mem_array[41573] = 16'hd233;
mem_array[41572] = 16'h3dfe;
mem_array[41575] = 16'hde96;
mem_array[41574] = 16'h3ed0;
mem_array[41577] = 16'hbb86;
mem_array[41576] = 16'hbef3;
mem_array[41579] = 16'h61fd;
mem_array[41578] = 16'h3dbf;
mem_array[41581] = 16'hf68d;
mem_array[41580] = 16'hbe85;
mem_array[41583] = 16'h0082;
mem_array[41582] = 16'h3b81;
mem_array[41585] = 16'h239d;
mem_array[41584] = 16'h3f71;
mem_array[41587] = 16'hbe59;
mem_array[41586] = 16'hbfb0;
mem_array[41589] = 16'h0320;
mem_array[41588] = 16'hbdb1;
mem_array[41591] = 16'hf6e9;
mem_array[41590] = 16'hbfcb;
mem_array[41593] = 16'h91a0;
mem_array[41592] = 16'h3de2;
mem_array[41595] = 16'h1497;
mem_array[41594] = 16'hbd14;
mem_array[41597] = 16'h89a8;
mem_array[41596] = 16'hbe8a;
mem_array[41599] = 16'h3fdf;
mem_array[41598] = 16'hbf90;
mem_array[41601] = 16'h3164;
mem_array[41600] = 16'h3d34;
mem_array[41603] = 16'heef6;
mem_array[41602] = 16'hbc6c;
mem_array[41605] = 16'h2daf;
mem_array[41604] = 16'hc012;
mem_array[41607] = 16'h611c;
mem_array[41606] = 16'hbe69;
mem_array[41609] = 16'h9e0f;
mem_array[41608] = 16'h3fa1;
mem_array[41611] = 16'hc507;
mem_array[41610] = 16'h3ec7;
mem_array[41613] = 16'h6774;
mem_array[41612] = 16'h3f5e;
mem_array[41615] = 16'h572f;
mem_array[41614] = 16'h3ed3;
mem_array[41617] = 16'h8657;
mem_array[41616] = 16'hbe35;
mem_array[41619] = 16'h2ab4;
mem_array[41618] = 16'hbebe;
mem_array[41621] = 16'hf019;
mem_array[41620] = 16'h3f78;
mem_array[41623] = 16'h85c9;
mem_array[41622] = 16'h3ea7;
mem_array[41625] = 16'h8dd5;
mem_array[41624] = 16'hbec1;
mem_array[41627] = 16'h8ed0;
mem_array[41626] = 16'hbe23;
mem_array[41629] = 16'hbd17;
mem_array[41628] = 16'hbf37;
mem_array[41631] = 16'h70c8;
mem_array[41630] = 16'hbfa3;
mem_array[41633] = 16'h72a1;
mem_array[41632] = 16'hbdbc;
mem_array[41635] = 16'hbebf;
mem_array[41634] = 16'h3ec5;
mem_array[41637] = 16'h743a;
mem_array[41636] = 16'h3dd8;
mem_array[41639] = 16'he314;
mem_array[41638] = 16'hbdbc;
mem_array[41641] = 16'h7568;
mem_array[41640] = 16'h3e9f;
mem_array[41643] = 16'h8b8f;
mem_array[41642] = 16'h3d3b;
mem_array[41645] = 16'hc19d;
mem_array[41644] = 16'h3f90;
mem_array[41647] = 16'he9cc;
mem_array[41646] = 16'hbf95;
mem_array[41649] = 16'h443d;
mem_array[41648] = 16'h3e4c;
mem_array[41651] = 16'hd3ea;
mem_array[41650] = 16'hbe80;
mem_array[41653] = 16'h5718;
mem_array[41652] = 16'h3f2f;
mem_array[41655] = 16'h5f04;
mem_array[41654] = 16'hbcce;
mem_array[41657] = 16'h78a5;
mem_array[41656] = 16'h3da9;
mem_array[41659] = 16'hcdaf;
mem_array[41658] = 16'hbf1a;
mem_array[41661] = 16'h5bf1;
mem_array[41660] = 16'hbd46;
mem_array[41663] = 16'h342f;
mem_array[41662] = 16'h3ce4;
mem_array[41665] = 16'hd809;
mem_array[41664] = 16'hbf11;
mem_array[41667] = 16'h0fcb;
mem_array[41666] = 16'h3e9e;
mem_array[41669] = 16'h8410;
mem_array[41668] = 16'h3f11;
mem_array[41671] = 16'h1bc4;
mem_array[41670] = 16'hbe1c;
mem_array[41673] = 16'hc496;
mem_array[41672] = 16'h3f18;
mem_array[41675] = 16'hc6c9;
mem_array[41674] = 16'hbe35;
mem_array[41677] = 16'h543f;
mem_array[41676] = 16'hbd46;
mem_array[41679] = 16'h2b83;
mem_array[41678] = 16'hbea6;
mem_array[41681] = 16'h3e7d;
mem_array[41680] = 16'h3f42;
mem_array[41683] = 16'h5ccd;
mem_array[41682] = 16'h3f00;
mem_array[41685] = 16'hd441;
mem_array[41684] = 16'hbecb;
mem_array[41687] = 16'hbca3;
mem_array[41686] = 16'hbe2f;
mem_array[41689] = 16'h9652;
mem_array[41688] = 16'hbea9;
mem_array[41691] = 16'h64df;
mem_array[41690] = 16'h3de4;
mem_array[41693] = 16'h690f;
mem_array[41692] = 16'h3e90;
mem_array[41695] = 16'h2ff2;
mem_array[41694] = 16'h3f34;
mem_array[41697] = 16'hb52a;
mem_array[41696] = 16'h3e55;
mem_array[41699] = 16'h83af;
mem_array[41698] = 16'hbf2b;
mem_array[41701] = 16'h5816;
mem_array[41700] = 16'h3f13;
mem_array[41703] = 16'hd7e3;
mem_array[41702] = 16'hbfa5;
mem_array[41705] = 16'h337a;
mem_array[41704] = 16'h3f01;
mem_array[41707] = 16'h9403;
mem_array[41706] = 16'hbfcd;
mem_array[41709] = 16'h98b2;
mem_array[41708] = 16'h3efa;
mem_array[41711] = 16'h57b1;
mem_array[41710] = 16'hbf17;
mem_array[41713] = 16'hc88f;
mem_array[41712] = 16'hbf1a;
mem_array[41715] = 16'h9481;
mem_array[41714] = 16'hbee9;
mem_array[41717] = 16'h1273;
mem_array[41716] = 16'h3db3;
mem_array[41719] = 16'h05c5;
mem_array[41718] = 16'h3f20;
mem_array[41721] = 16'hd500;
mem_array[41720] = 16'h3ac3;
mem_array[41723] = 16'hfc49;
mem_array[41722] = 16'hbc82;
mem_array[41725] = 16'h0fdf;
mem_array[41724] = 16'hbf5d;
mem_array[41727] = 16'haa40;
mem_array[41726] = 16'hbfc9;
mem_array[41729] = 16'he197;
mem_array[41728] = 16'h3f0d;
mem_array[41731] = 16'h0f65;
mem_array[41730] = 16'h3e94;
mem_array[41733] = 16'h47a5;
mem_array[41732] = 16'h3f68;
mem_array[41735] = 16'h8e67;
mem_array[41734] = 16'hbe9c;
mem_array[41737] = 16'hd3fa;
mem_array[41736] = 16'h3f2a;
mem_array[41739] = 16'ha158;
mem_array[41738] = 16'h3e5f;
mem_array[41741] = 16'hebdd;
mem_array[41740] = 16'h3ee6;
mem_array[41743] = 16'he76c;
mem_array[41742] = 16'h3e22;
mem_array[41745] = 16'hfaab;
mem_array[41744] = 16'hbef6;
mem_array[41747] = 16'h2446;
mem_array[41746] = 16'hbefb;
mem_array[41749] = 16'h83f4;
mem_array[41748] = 16'hbcfc;
mem_array[41751] = 16'hec97;
mem_array[41750] = 16'hbedb;
mem_array[41753] = 16'hec0b;
mem_array[41752] = 16'hbd3f;
mem_array[41755] = 16'he832;
mem_array[41754] = 16'hbd1a;
mem_array[41757] = 16'h4174;
mem_array[41756] = 16'hbeb6;
mem_array[41759] = 16'h6b3b;
mem_array[41758] = 16'hbf01;
mem_array[41761] = 16'hb9b5;
mem_array[41760] = 16'h3ef6;
mem_array[41763] = 16'h9bed;
mem_array[41762] = 16'h3de9;
mem_array[41765] = 16'hd4aa;
mem_array[41764] = 16'h3fae;
mem_array[41767] = 16'h7005;
mem_array[41766] = 16'hbe0e;
mem_array[41769] = 16'hb54b;
mem_array[41768] = 16'h3f00;
mem_array[41771] = 16'hb5b3;
mem_array[41770] = 16'hbf08;
mem_array[41773] = 16'h8b04;
mem_array[41772] = 16'h3cb1;
mem_array[41775] = 16'hf1bb;
mem_array[41774] = 16'hbeb4;
mem_array[41777] = 16'h3d58;
mem_array[41776] = 16'h3f40;
mem_array[41779] = 16'hb8fb;
mem_array[41778] = 16'h3ed5;
mem_array[41781] = 16'ha514;
mem_array[41780] = 16'hbd99;
mem_array[41783] = 16'h740f;
mem_array[41782] = 16'h3b99;
mem_array[41785] = 16'h9f07;
mem_array[41784] = 16'hbeb0;
mem_array[41787] = 16'h0086;
mem_array[41786] = 16'h3f8b;
mem_array[41789] = 16'h0e4a;
mem_array[41788] = 16'h3fba;
mem_array[41791] = 16'he7a0;
mem_array[41790] = 16'hbf23;
mem_array[41793] = 16'h6e09;
mem_array[41792] = 16'h400e;
mem_array[41795] = 16'h549e;
mem_array[41794] = 16'hbf8b;
mem_array[41797] = 16'h9ca6;
mem_array[41796] = 16'hbfa3;
mem_array[41799] = 16'hc9f4;
mem_array[41798] = 16'hbf64;
mem_array[41801] = 16'h386f;
mem_array[41800] = 16'hbf22;
mem_array[41803] = 16'h23b3;
mem_array[41802] = 16'h3eb5;
mem_array[41805] = 16'h1ec8;
mem_array[41804] = 16'hbcc4;
mem_array[41807] = 16'ha106;
mem_array[41806] = 16'hbeb6;
mem_array[41809] = 16'h8a51;
mem_array[41808] = 16'h3fa0;
mem_array[41811] = 16'hda02;
mem_array[41810] = 16'h3f21;
mem_array[41813] = 16'h2f5b;
mem_array[41812] = 16'h3f6f;
mem_array[41815] = 16'hec9a;
mem_array[41814] = 16'hbf17;
mem_array[41817] = 16'h13e1;
mem_array[41816] = 16'hbd03;
mem_array[41819] = 16'h6128;
mem_array[41818] = 16'hbe9b;
mem_array[41821] = 16'h82db;
mem_array[41820] = 16'hbd39;
mem_array[41823] = 16'h8ba2;
mem_array[41822] = 16'h3b65;
mem_array[41825] = 16'h01b2;
mem_array[41824] = 16'h3f7e;
mem_array[41827] = 16'h9869;
mem_array[41826] = 16'hbe1f;
mem_array[41829] = 16'h2472;
mem_array[41828] = 16'h3f60;
mem_array[41831] = 16'h2e48;
mem_array[41830] = 16'h3e8c;
mem_array[41833] = 16'h43eb;
mem_array[41832] = 16'h3e1a;
mem_array[41835] = 16'hb51d;
mem_array[41834] = 16'hbd9d;
mem_array[41837] = 16'h1ba4;
mem_array[41836] = 16'h3eaf;
mem_array[41839] = 16'h6d92;
mem_array[41838] = 16'h3e96;
mem_array[41841] = 16'hbc54;
mem_array[41840] = 16'h3c81;
mem_array[41843] = 16'h5964;
mem_array[41842] = 16'h3dab;
mem_array[41845] = 16'hf8e1;
mem_array[41844] = 16'hbf1b;
mem_array[41847] = 16'hc266;
mem_array[41846] = 16'h3f5a;
mem_array[41849] = 16'ha7c0;
mem_array[41848] = 16'h3f22;
mem_array[41851] = 16'h0001;
mem_array[41850] = 16'h3e8f;
mem_array[41853] = 16'hf94b;
mem_array[41852] = 16'h3c2b;
mem_array[41855] = 16'hd71a;
mem_array[41854] = 16'h3e2d;
mem_array[41857] = 16'h78f0;
mem_array[41856] = 16'hbe75;
mem_array[41859] = 16'h217b;
mem_array[41858] = 16'hbddc;
mem_array[41861] = 16'h180b;
mem_array[41860] = 16'h3f7c;
mem_array[41863] = 16'hfb2e;
mem_array[41862] = 16'hbf34;
mem_array[41865] = 16'hf29b;
mem_array[41864] = 16'h3c9f;
mem_array[41867] = 16'h61d9;
mem_array[41866] = 16'hbf18;
mem_array[41869] = 16'h0ed0;
mem_array[41868] = 16'h3f5c;
mem_array[41871] = 16'h3e14;
mem_array[41870] = 16'h3f0a;
mem_array[41873] = 16'hca4b;
mem_array[41872] = 16'hbe82;
mem_array[41875] = 16'hae32;
mem_array[41874] = 16'h3d4b;
mem_array[41877] = 16'hc5d8;
mem_array[41876] = 16'h3d0b;
mem_array[41879] = 16'hcbaa;
mem_array[41878] = 16'h3d89;
mem_array[41881] = 16'h5c02;
mem_array[41880] = 16'hbdd9;
mem_array[41883] = 16'he88a;
mem_array[41882] = 16'h3db8;
mem_array[41885] = 16'hd4ba;
mem_array[41884] = 16'h3f3d;
mem_array[41887] = 16'hba00;
mem_array[41886] = 16'hbbe8;
mem_array[41889] = 16'h314c;
mem_array[41888] = 16'hbd96;
mem_array[41891] = 16'hce17;
mem_array[41890] = 16'h3e41;
mem_array[41893] = 16'h4d02;
mem_array[41892] = 16'h3d25;
mem_array[41895] = 16'h72d1;
mem_array[41894] = 16'hbc07;
mem_array[41897] = 16'h2d97;
mem_array[41896] = 16'h3d03;
mem_array[41899] = 16'h952b;
mem_array[41898] = 16'h3e9b;
mem_array[41901] = 16'h14ff;
mem_array[41900] = 16'hbca7;
mem_array[41903] = 16'h2778;
mem_array[41902] = 16'h3d37;
mem_array[41905] = 16'ha203;
mem_array[41904] = 16'hbcda;
mem_array[41907] = 16'h19e6;
mem_array[41906] = 16'h3f58;
mem_array[41909] = 16'h44fe;
mem_array[41908] = 16'h3ef0;
mem_array[41911] = 16'haf16;
mem_array[41910] = 16'h3e8c;
mem_array[41913] = 16'h442a;
mem_array[41912] = 16'h3d95;
mem_array[41915] = 16'h792f;
mem_array[41914] = 16'hbbea;
mem_array[41917] = 16'hbc30;
mem_array[41916] = 16'hbe95;
mem_array[41919] = 16'h3148;
mem_array[41918] = 16'hbcbe;
mem_array[41921] = 16'h463c;
mem_array[41920] = 16'hbdf1;
mem_array[41923] = 16'h490e;
mem_array[41922] = 16'hbf01;
mem_array[41925] = 16'h27ef;
mem_array[41924] = 16'hbcc6;
mem_array[41927] = 16'h8331;
mem_array[41926] = 16'hbf69;
mem_array[41929] = 16'h9a64;
mem_array[41928] = 16'h3f63;
mem_array[41931] = 16'h0498;
mem_array[41930] = 16'h3cd9;
mem_array[41933] = 16'h5cc3;
mem_array[41932] = 16'h3f21;
mem_array[41935] = 16'hc375;
mem_array[41934] = 16'hbe84;
mem_array[41937] = 16'h3052;
mem_array[41936] = 16'h3b75;
mem_array[41939] = 16'hca4a;
mem_array[41938] = 16'hbd35;
mem_array[41941] = 16'h30b4;
mem_array[41940] = 16'h3ddf;
mem_array[41943] = 16'h5680;
mem_array[41942] = 16'hbd94;
mem_array[41945] = 16'hc924;
mem_array[41944] = 16'hbd20;
mem_array[41947] = 16'heff6;
mem_array[41946] = 16'hbc10;
mem_array[41949] = 16'hb4a1;
mem_array[41948] = 16'h3d5c;
mem_array[41951] = 16'h58d8;
mem_array[41950] = 16'hbcff;
mem_array[41953] = 16'h00e9;
mem_array[41952] = 16'h384f;
mem_array[41955] = 16'h084b;
mem_array[41954] = 16'hbb50;
mem_array[41957] = 16'hf4d1;
mem_array[41956] = 16'h3cbe;
mem_array[41959] = 16'h45df;
mem_array[41958] = 16'hbd85;
mem_array[41961] = 16'hb0da;
mem_array[41960] = 16'h3ce2;
mem_array[41963] = 16'hd474;
mem_array[41962] = 16'hbc1f;
mem_array[41965] = 16'hdafd;
mem_array[41964] = 16'hbd62;
mem_array[41967] = 16'h44ca;
mem_array[41966] = 16'hbda0;
mem_array[41969] = 16'ha3b7;
mem_array[41968] = 16'hbd34;
mem_array[41971] = 16'hc657;
mem_array[41970] = 16'h3c3e;
mem_array[41973] = 16'h7816;
mem_array[41972] = 16'hbce8;
mem_array[41975] = 16'h34c5;
mem_array[41974] = 16'h3c9a;
mem_array[41977] = 16'h14d5;
mem_array[41976] = 16'h3b1e;
mem_array[41979] = 16'h35c7;
mem_array[41978] = 16'h3be0;
mem_array[41981] = 16'hd201;
mem_array[41980] = 16'h3db5;
mem_array[41983] = 16'h911b;
mem_array[41982] = 16'h3d66;
mem_array[41985] = 16'h8d45;
mem_array[41984] = 16'h3c86;
mem_array[41987] = 16'hf072;
mem_array[41986] = 16'h3d81;
mem_array[41989] = 16'h8723;
mem_array[41988] = 16'hbbea;
mem_array[41991] = 16'h4ddc;
mem_array[41990] = 16'h3b11;
mem_array[41993] = 16'hc889;
mem_array[41992] = 16'hbc6c;
mem_array[41995] = 16'h4964;
mem_array[41994] = 16'h3d6d;
mem_array[41997] = 16'h682f;
mem_array[41996] = 16'hbbdd;
mem_array[41999] = 16'h9c83;
mem_array[41998] = 16'h3d91;
mem_array[42001] = 16'h62d1;
mem_array[42000] = 16'h3ca3;
mem_array[42003] = 16'hb996;
mem_array[42002] = 16'h3baa;
mem_array[42005] = 16'hdf6d;
mem_array[42004] = 16'hbc7d;
mem_array[42007] = 16'ha428;
mem_array[42006] = 16'h3d1f;
mem_array[42009] = 16'hcff8;
mem_array[42008] = 16'h3c80;
mem_array[42011] = 16'hd121;
mem_array[42010] = 16'h3d2d;
mem_array[42013] = 16'h4fe8;
mem_array[42012] = 16'h3ccd;
mem_array[42015] = 16'h5c33;
mem_array[42014] = 16'h3c75;
mem_array[42017] = 16'h58a4;
mem_array[42016] = 16'hbc51;
mem_array[42019] = 16'hfd12;
mem_array[42018] = 16'h3c0e;
mem_array[42021] = 16'hd567;
mem_array[42020] = 16'h3ccd;
mem_array[42023] = 16'hdbb5;
mem_array[42022] = 16'hbcc9;
mem_array[42025] = 16'he35c;
mem_array[42024] = 16'hbd6c;
mem_array[42027] = 16'h5cc4;
mem_array[42026] = 16'h3d9d;
mem_array[42029] = 16'h1687;
mem_array[42028] = 16'h3bd7;
mem_array[42031] = 16'h7c58;
mem_array[42030] = 16'hbca6;
mem_array[42033] = 16'hd832;
mem_array[42032] = 16'hbd6f;
mem_array[42035] = 16'h600f;
mem_array[42034] = 16'h3c73;
mem_array[42037] = 16'h7bff;
mem_array[42036] = 16'h3d24;
mem_array[42039] = 16'h8503;
mem_array[42038] = 16'hbcee;
mem_array[42041] = 16'h3513;
mem_array[42040] = 16'hbdc0;
mem_array[42043] = 16'ha93d;
mem_array[42042] = 16'hbbeb;
mem_array[42045] = 16'ha08d;
mem_array[42044] = 16'hbcf7;
mem_array[42047] = 16'h2cc4;
mem_array[42046] = 16'h3d39;
mem_array[42049] = 16'h036d;
mem_array[42048] = 16'hbd83;
mem_array[42051] = 16'h6540;
mem_array[42050] = 16'hbb91;
mem_array[42053] = 16'haaa1;
mem_array[42052] = 16'h3d0d;
mem_array[42055] = 16'hf52d;
mem_array[42054] = 16'hbd38;
mem_array[42057] = 16'h6470;
mem_array[42056] = 16'h3dac;
mem_array[42059] = 16'h69e2;
mem_array[42058] = 16'hbcb0;
mem_array[42061] = 16'hec08;
mem_array[42060] = 16'h3d2d;
mem_array[42063] = 16'haa35;
mem_array[42062] = 16'h3c91;
mem_array[42065] = 16'h47cf;
mem_array[42064] = 16'h3b0e;
mem_array[42067] = 16'h2151;
mem_array[42066] = 16'hbc2a;
mem_array[42069] = 16'ha99b;
mem_array[42068] = 16'hbb7e;
mem_array[42071] = 16'h6379;
mem_array[42070] = 16'h3cf1;
mem_array[42073] = 16'hafe2;
mem_array[42072] = 16'h3d19;
mem_array[42075] = 16'hf03b;
mem_array[42074] = 16'hbbe9;
mem_array[42077] = 16'h2564;
mem_array[42076] = 16'hbc4c;
mem_array[42079] = 16'h5df8;
mem_array[42078] = 16'hbc38;
mem_array[42081] = 16'h2ce6;
mem_array[42080] = 16'hba09;
mem_array[42083] = 16'h31da;
mem_array[42082] = 16'hbd87;
mem_array[42085] = 16'h95cc;
mem_array[42084] = 16'h3d8f;
mem_array[42087] = 16'h090c;
mem_array[42086] = 16'h3d78;
mem_array[42089] = 16'h470f;
mem_array[42088] = 16'h3cc1;
mem_array[42091] = 16'h8d02;
mem_array[42090] = 16'h3d92;
mem_array[42093] = 16'h35bd;
mem_array[42092] = 16'hbd4d;
mem_array[42095] = 16'h26ba;
mem_array[42094] = 16'h3d80;
mem_array[42097] = 16'h281a;
mem_array[42096] = 16'hbd00;
mem_array[42099] = 16'h551f;
mem_array[42098] = 16'hbcf8;
mem_array[42101] = 16'h625f;
mem_array[42100] = 16'hbc31;
mem_array[42103] = 16'hf997;
mem_array[42102] = 16'h3d3c;
mem_array[42105] = 16'h89e8;
mem_array[42104] = 16'h3dae;
mem_array[42107] = 16'h4422;
mem_array[42106] = 16'h3dc5;
mem_array[42109] = 16'h41b4;
mem_array[42108] = 16'h3da9;
mem_array[42111] = 16'h1420;
mem_array[42110] = 16'h3d0a;
mem_array[42113] = 16'hbb93;
mem_array[42112] = 16'hbcb0;
mem_array[42115] = 16'h154a;
mem_array[42114] = 16'hbd99;
mem_array[42117] = 16'hd46c;
mem_array[42116] = 16'hbcc4;
mem_array[42119] = 16'h148a;
mem_array[42118] = 16'h3baa;
mem_array[42121] = 16'h78e7;
mem_array[42120] = 16'hbcdc;
mem_array[42123] = 16'h0195;
mem_array[42122] = 16'h3e1b;
mem_array[42125] = 16'hdd01;
mem_array[42124] = 16'hbd56;
mem_array[42127] = 16'he40e;
mem_array[42126] = 16'hbd6e;
mem_array[42129] = 16'h1605;
mem_array[42128] = 16'hbcf4;
mem_array[42131] = 16'he45a;
mem_array[42130] = 16'hbe12;
mem_array[42133] = 16'h3a69;
mem_array[42132] = 16'h3ea6;
mem_array[42135] = 16'h184a;
mem_array[42134] = 16'hbd12;
mem_array[42137] = 16'h3023;
mem_array[42136] = 16'hbcab;
mem_array[42139] = 16'he10d;
mem_array[42138] = 16'h3d64;
mem_array[42141] = 16'h0f97;
mem_array[42140] = 16'h3cc5;
mem_array[42143] = 16'h5ff4;
mem_array[42142] = 16'h3cad;
mem_array[42145] = 16'h6c16;
mem_array[42144] = 16'hbd99;
mem_array[42147] = 16'he604;
mem_array[42146] = 16'h3dd8;
mem_array[42149] = 16'he1f8;
mem_array[42148] = 16'hbdd8;
mem_array[42151] = 16'hec41;
mem_array[42150] = 16'h3bd8;
mem_array[42153] = 16'h019b;
mem_array[42152] = 16'hbda6;
mem_array[42155] = 16'hdec1;
mem_array[42154] = 16'h3d48;
mem_array[42157] = 16'hef00;
mem_array[42156] = 16'h3f13;
mem_array[42159] = 16'hd3da;
mem_array[42158] = 16'hbeba;
mem_array[42161] = 16'haa72;
mem_array[42160] = 16'h3b86;
mem_array[42163] = 16'h1a82;
mem_array[42162] = 16'h3e17;
mem_array[42165] = 16'h3088;
mem_array[42164] = 16'h3cea;
mem_array[42167] = 16'h833e;
mem_array[42166] = 16'hbf4f;
mem_array[42169] = 16'h132e;
mem_array[42168] = 16'h3e95;
mem_array[42171] = 16'h5f9c;
mem_array[42170] = 16'hbdde;
mem_array[42173] = 16'hff7c;
mem_array[42172] = 16'h3ec8;
mem_array[42175] = 16'hb347;
mem_array[42174] = 16'h3d64;
mem_array[42177] = 16'h00ce;
mem_array[42176] = 16'hbca9;
mem_array[42179] = 16'hdb2c;
mem_array[42178] = 16'hbcaa;
mem_array[42181] = 16'h9c7e;
mem_array[42180] = 16'h3dfa;
mem_array[42183] = 16'hdd36;
mem_array[42182] = 16'hbc80;
mem_array[42185] = 16'h3d08;
mem_array[42184] = 16'h3df4;
mem_array[42187] = 16'h0de7;
mem_array[42186] = 16'h3d50;
mem_array[42189] = 16'h7db1;
mem_array[42188] = 16'h3f93;
mem_array[42191] = 16'hac85;
mem_array[42190] = 16'h3ebf;
mem_array[42193] = 16'h1abe;
mem_array[42192] = 16'h3c03;
mem_array[42195] = 16'h9860;
mem_array[42194] = 16'hbe9f;
mem_array[42197] = 16'hf308;
mem_array[42196] = 16'hbe2f;
mem_array[42199] = 16'h9dc3;
mem_array[42198] = 16'hbcb4;
mem_array[42201] = 16'h13e0;
mem_array[42200] = 16'hbc98;
mem_array[42203] = 16'h9c41;
mem_array[42202] = 16'hbbfc;
mem_array[42205] = 16'hceab;
mem_array[42204] = 16'h3c15;
mem_array[42207] = 16'ha05f;
mem_array[42206] = 16'hbddb;
mem_array[42209] = 16'h6f63;
mem_array[42208] = 16'h3ca9;
mem_array[42211] = 16'hd89b;
mem_array[42210] = 16'hbe9f;
mem_array[42213] = 16'h952b;
mem_array[42212] = 16'hbe49;
mem_array[42215] = 16'h95bf;
mem_array[42214] = 16'hbcb3;
mem_array[42217] = 16'h5e00;
mem_array[42216] = 16'h3e64;
mem_array[42219] = 16'hd123;
mem_array[42218] = 16'h3d47;
mem_array[42221] = 16'h6770;
mem_array[42220] = 16'hbd0f;
mem_array[42223] = 16'h7f39;
mem_array[42222] = 16'hbed8;
mem_array[42225] = 16'hae0f;
mem_array[42224] = 16'h3dd7;
mem_array[42227] = 16'ha677;
mem_array[42226] = 16'hbd7f;
mem_array[42229] = 16'hd0b5;
mem_array[42228] = 16'hbddb;
mem_array[42231] = 16'h6f5b;
mem_array[42230] = 16'h3f42;
mem_array[42233] = 16'h4bc6;
mem_array[42232] = 16'hbf31;
mem_array[42235] = 16'hf3fb;
mem_array[42234] = 16'h3e03;
mem_array[42237] = 16'h6a9f;
mem_array[42236] = 16'hbd1c;
mem_array[42239] = 16'hb568;
mem_array[42238] = 16'hbe0b;
mem_array[42241] = 16'h4a7c;
mem_array[42240] = 16'hbf19;
mem_array[42243] = 16'ha6e0;
mem_array[42242] = 16'h3f6f;
mem_array[42245] = 16'h25ef;
mem_array[42244] = 16'hbee6;
mem_array[42247] = 16'h01c9;
mem_array[42246] = 16'hbe9f;
mem_array[42249] = 16'h54d9;
mem_array[42248] = 16'h3f71;
mem_array[42251] = 16'h518a;
mem_array[42250] = 16'h3d81;
mem_array[42253] = 16'h690f;
mem_array[42252] = 16'h3fdb;
mem_array[42255] = 16'h8bde;
mem_array[42254] = 16'hbe98;
mem_array[42257] = 16'hc528;
mem_array[42256] = 16'hbd49;
mem_array[42259] = 16'hb1ef;
mem_array[42258] = 16'h3c45;
mem_array[42261] = 16'haa93;
mem_array[42260] = 16'hb985;
mem_array[42263] = 16'h4604;
mem_array[42262] = 16'h3acc;
mem_array[42265] = 16'he12e;
mem_array[42264] = 16'hbe53;
mem_array[42267] = 16'hc3f4;
mem_array[42266] = 16'hbe50;
mem_array[42269] = 16'h484d;
mem_array[42268] = 16'hbec9;
mem_array[42271] = 16'he9fd;
mem_array[42270] = 16'h3f1c;
mem_array[42273] = 16'h421c;
mem_array[42272] = 16'hbf5e;
mem_array[42275] = 16'hdb9d;
mem_array[42274] = 16'hbed2;
mem_array[42277] = 16'h093a;
mem_array[42276] = 16'hbef1;
mem_array[42279] = 16'hf8c3;
mem_array[42278] = 16'h3b36;
mem_array[42281] = 16'h6225;
mem_array[42280] = 16'hbf36;
mem_array[42283] = 16'h88c8;
mem_array[42282] = 16'h3eef;
mem_array[42285] = 16'h5e26;
mem_array[42284] = 16'h3d14;
mem_array[42287] = 16'h8431;
mem_array[42286] = 16'h3e21;
mem_array[42289] = 16'h97f9;
mem_array[42288] = 16'h3f02;
mem_array[42291] = 16'hd108;
mem_array[42290] = 16'hbda4;
mem_array[42293] = 16'h5ece;
mem_array[42292] = 16'hbea4;
mem_array[42295] = 16'h3fdc;
mem_array[42294] = 16'hbe12;
mem_array[42297] = 16'h8868;
mem_array[42296] = 16'hbde7;
mem_array[42299] = 16'h6d28;
mem_array[42298] = 16'h3e26;
mem_array[42301] = 16'hd765;
mem_array[42300] = 16'hbe81;
mem_array[42303] = 16'h47ad;
mem_array[42302] = 16'h3e92;
mem_array[42305] = 16'h9539;
mem_array[42304] = 16'hbf7f;
mem_array[42307] = 16'h9d77;
mem_array[42306] = 16'hbdec;
mem_array[42309] = 16'heb07;
mem_array[42308] = 16'h3f3e;
mem_array[42311] = 16'h4bd7;
mem_array[42310] = 16'hbe56;
mem_array[42313] = 16'h75f3;
mem_array[42312] = 16'h3f3e;
mem_array[42315] = 16'h32b5;
mem_array[42314] = 16'hbe53;
mem_array[42317] = 16'h1709;
mem_array[42316] = 16'hbe23;
mem_array[42319] = 16'hdd69;
mem_array[42318] = 16'hbe0d;
mem_array[42321] = 16'h0cda;
mem_array[42320] = 16'h3dbd;
mem_array[42323] = 16'hd4fb;
mem_array[42322] = 16'hbdb0;
mem_array[42325] = 16'h18ac;
mem_array[42324] = 16'hbfac;
mem_array[42327] = 16'h1add;
mem_array[42326] = 16'hbf94;
mem_array[42329] = 16'h7f63;
mem_array[42328] = 16'hbe5b;
mem_array[42331] = 16'h54bd;
mem_array[42330] = 16'hbe6a;
mem_array[42333] = 16'hb402;
mem_array[42332] = 16'hbf9d;
mem_array[42335] = 16'h87ec;
mem_array[42334] = 16'hbf3e;
mem_array[42337] = 16'hd47b;
mem_array[42336] = 16'hbe96;
mem_array[42339] = 16'hdf3b;
mem_array[42338] = 16'h3d8c;
mem_array[42341] = 16'h22ba;
mem_array[42340] = 16'hbf72;
mem_array[42343] = 16'h6e30;
mem_array[42342] = 16'h3f09;
mem_array[42345] = 16'h3a4a;
mem_array[42344] = 16'hbc93;
mem_array[42347] = 16'h377e;
mem_array[42346] = 16'h3f14;
mem_array[42349] = 16'h5548;
mem_array[42348] = 16'h3e57;
mem_array[42351] = 16'hfc14;
mem_array[42350] = 16'hbf7a;
mem_array[42353] = 16'h10cf;
mem_array[42352] = 16'h3e02;
mem_array[42355] = 16'h2875;
mem_array[42354] = 16'hbe12;
mem_array[42357] = 16'h9bab;
mem_array[42356] = 16'hbe82;
mem_array[42359] = 16'hff04;
mem_array[42358] = 16'h3e09;
mem_array[42361] = 16'hbe1f;
mem_array[42360] = 16'hbe97;
mem_array[42363] = 16'haa19;
mem_array[42362] = 16'h3eb8;
mem_array[42365] = 16'h4060;
mem_array[42364] = 16'hbe43;
mem_array[42367] = 16'hafaa;
mem_array[42366] = 16'hbed8;
mem_array[42369] = 16'ha9f7;
mem_array[42368] = 16'h3e02;
mem_array[42371] = 16'h3588;
mem_array[42370] = 16'hbe95;
mem_array[42373] = 16'ha8bb;
mem_array[42372] = 16'h3edb;
mem_array[42375] = 16'ha839;
mem_array[42374] = 16'h3d12;
mem_array[42377] = 16'h41d9;
mem_array[42376] = 16'hbf42;
mem_array[42379] = 16'h4233;
mem_array[42378] = 16'hbe40;
mem_array[42381] = 16'hded4;
mem_array[42380] = 16'h3d6f;
mem_array[42383] = 16'hef0f;
mem_array[42382] = 16'hbd20;
mem_array[42385] = 16'hdde9;
mem_array[42384] = 16'hbfc1;
mem_array[42387] = 16'h61c1;
mem_array[42386] = 16'hbf5f;
mem_array[42389] = 16'hfd0b;
mem_array[42388] = 16'h3efe;
mem_array[42391] = 16'hde67;
mem_array[42390] = 16'hbf02;
mem_array[42393] = 16'hdabc;
mem_array[42392] = 16'hbfac;
mem_array[42395] = 16'h98f7;
mem_array[42394] = 16'hbf0a;
mem_array[42397] = 16'h2d65;
mem_array[42396] = 16'hbf48;
mem_array[42399] = 16'h7772;
mem_array[42398] = 16'h3e70;
mem_array[42401] = 16'hb326;
mem_array[42400] = 16'hbf43;
mem_array[42403] = 16'h619a;
mem_array[42402] = 16'h3f0b;
mem_array[42405] = 16'h71db;
mem_array[42404] = 16'hbd09;
mem_array[42407] = 16'hc8b9;
mem_array[42406] = 16'h3f72;
mem_array[42409] = 16'h6688;
mem_array[42408] = 16'h3ed5;
mem_array[42411] = 16'h201a;
mem_array[42410] = 16'hbeac;
mem_array[42413] = 16'hce68;
mem_array[42412] = 16'h3f2a;
mem_array[42415] = 16'h53f4;
mem_array[42414] = 16'h3d89;
mem_array[42417] = 16'h2881;
mem_array[42416] = 16'hbe99;
mem_array[42419] = 16'h7548;
mem_array[42418] = 16'h3dcc;
mem_array[42421] = 16'hc162;
mem_array[42420] = 16'hbce8;
mem_array[42423] = 16'hfbae;
mem_array[42422] = 16'h3e85;
mem_array[42425] = 16'h01ca;
mem_array[42424] = 16'hbcae;
mem_array[42427] = 16'h8193;
mem_array[42426] = 16'hbe65;
mem_array[42429] = 16'ha8f0;
mem_array[42428] = 16'h3eec;
mem_array[42431] = 16'hb3e4;
mem_array[42430] = 16'hbf24;
mem_array[42433] = 16'h981f;
mem_array[42432] = 16'h3f20;
mem_array[42435] = 16'h1be2;
mem_array[42434] = 16'h3e6f;
mem_array[42437] = 16'h389c;
mem_array[42436] = 16'hbf13;
mem_array[42439] = 16'h5cbe;
mem_array[42438] = 16'hbeac;
mem_array[42441] = 16'h21f4;
mem_array[42440] = 16'hbd19;
mem_array[42443] = 16'h40b8;
mem_array[42442] = 16'hbd8a;
mem_array[42445] = 16'hc305;
mem_array[42444] = 16'hbee6;
mem_array[42447] = 16'h9a27;
mem_array[42446] = 16'hbf6a;
mem_array[42449] = 16'h7bde;
mem_array[42448] = 16'h3f42;
mem_array[42451] = 16'h0c8e;
mem_array[42450] = 16'hbedf;
mem_array[42453] = 16'h85d0;
mem_array[42452] = 16'hbf82;
mem_array[42455] = 16'h73d4;
mem_array[42454] = 16'hbf14;
mem_array[42457] = 16'h1937;
mem_array[42456] = 16'hbeb7;
mem_array[42459] = 16'h1426;
mem_array[42458] = 16'h3f36;
mem_array[42461] = 16'h4655;
mem_array[42460] = 16'hbf10;
mem_array[42463] = 16'h3897;
mem_array[42462] = 16'h3f6c;
mem_array[42465] = 16'ha5a9;
mem_array[42464] = 16'h3c04;
mem_array[42467] = 16'h2722;
mem_array[42466] = 16'h3f1d;
mem_array[42469] = 16'h1453;
mem_array[42468] = 16'h3e98;
mem_array[42471] = 16'h8056;
mem_array[42470] = 16'h3e4a;
mem_array[42473] = 16'h64d1;
mem_array[42472] = 16'h3f1f;
mem_array[42475] = 16'hae4a;
mem_array[42474] = 16'hbcea;
mem_array[42477] = 16'he20d;
mem_array[42476] = 16'hbee4;
mem_array[42479] = 16'h81c2;
mem_array[42478] = 16'hbf61;
mem_array[42481] = 16'h244c;
mem_array[42480] = 16'h3f03;
mem_array[42483] = 16'h58df;
mem_array[42482] = 16'h3e09;
mem_array[42485] = 16'h0393;
mem_array[42484] = 16'h3eea;
mem_array[42487] = 16'ha40b;
mem_array[42486] = 16'hbf54;
mem_array[42489] = 16'h9682;
mem_array[42488] = 16'h3f0c;
mem_array[42491] = 16'h3273;
mem_array[42490] = 16'hbeaa;
mem_array[42493] = 16'h09df;
mem_array[42492] = 16'h3f41;
mem_array[42495] = 16'h3f19;
mem_array[42494] = 16'hbf5a;
mem_array[42497] = 16'h8d84;
mem_array[42496] = 16'hbf09;
mem_array[42499] = 16'h035c;
mem_array[42498] = 16'hbde8;
mem_array[42501] = 16'hd008;
mem_array[42500] = 16'hbd97;
mem_array[42503] = 16'hcc32;
mem_array[42502] = 16'hbc01;
mem_array[42505] = 16'h9512;
mem_array[42504] = 16'hbcae;
mem_array[42507] = 16'h54b7;
mem_array[42506] = 16'hbfac;
mem_array[42509] = 16'hf9ea;
mem_array[42508] = 16'h3f1a;
mem_array[42511] = 16'h23b1;
mem_array[42510] = 16'h3dad;
mem_array[42513] = 16'hecbe;
mem_array[42512] = 16'hbe71;
mem_array[42515] = 16'hd7ae;
mem_array[42514] = 16'hbed0;
mem_array[42517] = 16'hd6df;
mem_array[42516] = 16'hbd96;
mem_array[42519] = 16'h58de;
mem_array[42518] = 16'h3e2d;
mem_array[42521] = 16'h8225;
mem_array[42520] = 16'hbec9;
mem_array[42523] = 16'h46b0;
mem_array[42522] = 16'h3f07;
mem_array[42525] = 16'hc13d;
mem_array[42524] = 16'hbcbc;
mem_array[42527] = 16'h1188;
mem_array[42526] = 16'h3d7b;
mem_array[42529] = 16'h0344;
mem_array[42528] = 16'h3ef8;
mem_array[42531] = 16'h3037;
mem_array[42530] = 16'h3eac;
mem_array[42533] = 16'hac77;
mem_array[42532] = 16'h3ef4;
mem_array[42535] = 16'h3b40;
mem_array[42534] = 16'hbebd;
mem_array[42537] = 16'hf8e6;
mem_array[42536] = 16'hbf35;
mem_array[42539] = 16'h152e;
mem_array[42538] = 16'hbf39;
mem_array[42541] = 16'h7cf1;
mem_array[42540] = 16'h3e5c;
mem_array[42543] = 16'h045a;
mem_array[42542] = 16'h3e92;
mem_array[42545] = 16'h5c44;
mem_array[42544] = 16'h3e02;
mem_array[42547] = 16'hfd71;
mem_array[42546] = 16'hbf83;
mem_array[42549] = 16'h081c;
mem_array[42548] = 16'h3d51;
mem_array[42551] = 16'hc08a;
mem_array[42550] = 16'h3de9;
mem_array[42553] = 16'hd92e;
mem_array[42552] = 16'hbeb4;
mem_array[42555] = 16'h9396;
mem_array[42554] = 16'hbfd9;
mem_array[42557] = 16'h5053;
mem_array[42556] = 16'hbfc0;
mem_array[42559] = 16'hbaa3;
mem_array[42558] = 16'hbe0a;
mem_array[42561] = 16'h5ac8;
mem_array[42560] = 16'h3d7d;
mem_array[42563] = 16'h44ac;
mem_array[42562] = 16'hbc71;
mem_array[42565] = 16'h9af7;
mem_array[42564] = 16'hbfe7;
mem_array[42567] = 16'hc2ab;
mem_array[42566] = 16'hbfae;
mem_array[42569] = 16'h58c0;
mem_array[42568] = 16'hbeb5;
mem_array[42571] = 16'hc984;
mem_array[42570] = 16'hbe22;
mem_array[42573] = 16'hd296;
mem_array[42572] = 16'hbe0e;
mem_array[42575] = 16'h0456;
mem_array[42574] = 16'hbecf;
mem_array[42577] = 16'h0fcb;
mem_array[42576] = 16'h3db4;
mem_array[42579] = 16'h781f;
mem_array[42578] = 16'hbf93;
mem_array[42581] = 16'h25bb;
mem_array[42580] = 16'hbdbd;
mem_array[42583] = 16'h23f0;
mem_array[42582] = 16'h3f32;
mem_array[42585] = 16'hb9d0;
mem_array[42584] = 16'hbd1a;
mem_array[42587] = 16'hf4af;
mem_array[42586] = 16'h3e60;
mem_array[42589] = 16'h1cfa;
mem_array[42588] = 16'h3e11;
mem_array[42591] = 16'hab1c;
mem_array[42590] = 16'h3e7b;
mem_array[42593] = 16'he529;
mem_array[42592] = 16'h3ef5;
mem_array[42595] = 16'h3c59;
mem_array[42594] = 16'hbde6;
mem_array[42597] = 16'h2a8c;
mem_array[42596] = 16'hbf19;
mem_array[42599] = 16'h7246;
mem_array[42598] = 16'hbf78;
mem_array[42601] = 16'h5291;
mem_array[42600] = 16'hbcb6;
mem_array[42603] = 16'hd3cf;
mem_array[42602] = 16'h3e82;
mem_array[42605] = 16'h6222;
mem_array[42604] = 16'hbd07;
mem_array[42607] = 16'had12;
mem_array[42606] = 16'hbf9a;
mem_array[42609] = 16'hdf9a;
mem_array[42608] = 16'h3d6a;
mem_array[42611] = 16'h63d8;
mem_array[42610] = 16'h3e33;
mem_array[42613] = 16'h9f23;
mem_array[42612] = 16'h3efd;
mem_array[42615] = 16'h59b5;
mem_array[42614] = 16'hbf0e;
mem_array[42617] = 16'h9515;
mem_array[42616] = 16'hbf78;
mem_array[42619] = 16'ha2ba;
mem_array[42618] = 16'hc00d;
mem_array[42621] = 16'h2a92;
mem_array[42620] = 16'h3d8f;
mem_array[42623] = 16'h5aee;
mem_array[42622] = 16'h3cc2;
mem_array[42625] = 16'h453c;
mem_array[42624] = 16'hbf84;
mem_array[42627] = 16'ha1f7;
mem_array[42626] = 16'hbfa2;
mem_array[42629] = 16'h73ec;
mem_array[42628] = 16'hbf77;
mem_array[42631] = 16'h82c2;
mem_array[42630] = 16'hbe40;
mem_array[42633] = 16'h4a9a;
mem_array[42632] = 16'hbf77;
mem_array[42635] = 16'h32d6;
mem_array[42634] = 16'hbe71;
mem_array[42637] = 16'h541b;
mem_array[42636] = 16'hbec7;
mem_array[42639] = 16'hfdc1;
mem_array[42638] = 16'hbeac;
mem_array[42641] = 16'h33e2;
mem_array[42640] = 16'hbe2b;
mem_array[42643] = 16'hdb30;
mem_array[42642] = 16'h3ef2;
mem_array[42645] = 16'h9bcc;
mem_array[42644] = 16'h3bff;
mem_array[42647] = 16'h7da9;
mem_array[42646] = 16'h3ec4;
mem_array[42649] = 16'hcd38;
mem_array[42648] = 16'h3e6d;
mem_array[42651] = 16'heb92;
mem_array[42650] = 16'hbe0c;
mem_array[42653] = 16'h6a3d;
mem_array[42652] = 16'h3ec0;
mem_array[42655] = 16'he1ea;
mem_array[42654] = 16'h3e7e;
mem_array[42657] = 16'h8b40;
mem_array[42656] = 16'hbe98;
mem_array[42659] = 16'h3800;
mem_array[42658] = 16'hbf52;
mem_array[42661] = 16'h13bc;
mem_array[42660] = 16'h3e94;
mem_array[42663] = 16'hf6a1;
mem_array[42662] = 16'h3e9a;
mem_array[42665] = 16'h0cd8;
mem_array[42664] = 16'h3de0;
mem_array[42667] = 16'hae37;
mem_array[42666] = 16'hbfaf;
mem_array[42669] = 16'h8387;
mem_array[42668] = 16'h3ece;
mem_array[42671] = 16'hc83a;
mem_array[42670] = 16'h3dd2;
mem_array[42673] = 16'h1553;
mem_array[42672] = 16'h3dcb;
mem_array[42675] = 16'ha721;
mem_array[42674] = 16'h3daa;
mem_array[42677] = 16'haa5c;
mem_array[42676] = 16'h3ebc;
mem_array[42679] = 16'hda39;
mem_array[42678] = 16'hbff6;
mem_array[42681] = 16'h6ff5;
mem_array[42680] = 16'h3d8b;
mem_array[42683] = 16'h2520;
mem_array[42682] = 16'h3d10;
mem_array[42685] = 16'h7586;
mem_array[42684] = 16'hbfb2;
mem_array[42687] = 16'hd6c3;
mem_array[42686] = 16'hbf7d;
mem_array[42689] = 16'h0e09;
mem_array[42688] = 16'hbeff;
mem_array[42691] = 16'h3b6f;
mem_array[42690] = 16'hbeaa;
mem_array[42693] = 16'hb63a;
mem_array[42692] = 16'hbf7c;
mem_array[42695] = 16'h5b76;
mem_array[42694] = 16'h3d23;
mem_array[42697] = 16'habff;
mem_array[42696] = 16'hbe38;
mem_array[42699] = 16'h18b2;
mem_array[42698] = 16'hbea9;
mem_array[42701] = 16'h9ccf;
mem_array[42700] = 16'hbec0;
mem_array[42703] = 16'hdc07;
mem_array[42702] = 16'h3e8a;
mem_array[42705] = 16'h3700;
mem_array[42704] = 16'h3e80;
mem_array[42707] = 16'hbb5b;
mem_array[42706] = 16'h3e20;
mem_array[42709] = 16'h3622;
mem_array[42708] = 16'hbd4c;
mem_array[42711] = 16'h7128;
mem_array[42710] = 16'h3cc7;
mem_array[42713] = 16'h4ed4;
mem_array[42712] = 16'h3ea0;
mem_array[42715] = 16'h625a;
mem_array[42714] = 16'h3c97;
mem_array[42717] = 16'h01c9;
mem_array[42716] = 16'h3d06;
mem_array[42719] = 16'hfaf4;
mem_array[42718] = 16'hbf41;
mem_array[42721] = 16'h58a3;
mem_array[42720] = 16'h3e3e;
mem_array[42723] = 16'h69f1;
mem_array[42722] = 16'h3e7b;
mem_array[42725] = 16'h2ec2;
mem_array[42724] = 16'h3ee9;
mem_array[42727] = 16'hcfe6;
mem_array[42726] = 16'hbf62;
mem_array[42729] = 16'h8c42;
mem_array[42728] = 16'h3e0a;
mem_array[42731] = 16'h6abc;
mem_array[42730] = 16'h3f1e;
mem_array[42733] = 16'h9f17;
mem_array[42732] = 16'hbe72;
mem_array[42735] = 16'hb946;
mem_array[42734] = 16'h3d7c;
mem_array[42737] = 16'h37c2;
mem_array[42736] = 16'h3e8b;
mem_array[42739] = 16'hd802;
mem_array[42738] = 16'hbfe8;
mem_array[42741] = 16'ha30d;
mem_array[42740] = 16'hbdb1;
mem_array[42743] = 16'h44fc;
mem_array[42742] = 16'h3c84;
mem_array[42745] = 16'h2126;
mem_array[42744] = 16'hc007;
mem_array[42747] = 16'hed2b;
mem_array[42746] = 16'hbf5a;
mem_array[42749] = 16'hcb93;
mem_array[42748] = 16'h3ee6;
mem_array[42751] = 16'h6e0e;
mem_array[42750] = 16'hbeb6;
mem_array[42753] = 16'h5b55;
mem_array[42752] = 16'hbfa8;
mem_array[42755] = 16'h5124;
mem_array[42754] = 16'hbce0;
mem_array[42757] = 16'h88ad;
mem_array[42756] = 16'hbca8;
mem_array[42759] = 16'h4493;
mem_array[42758] = 16'hbe93;
mem_array[42761] = 16'hb051;
mem_array[42760] = 16'hbe8e;
mem_array[42763] = 16'h93b8;
mem_array[42762] = 16'h3e1b;
mem_array[42765] = 16'hcd10;
mem_array[42764] = 16'hbe2b;
mem_array[42767] = 16'hc7ed;
mem_array[42766] = 16'hbe9e;
mem_array[42769] = 16'h0df7;
mem_array[42768] = 16'h3e4e;
mem_array[42771] = 16'h633a;
mem_array[42770] = 16'h3e98;
mem_array[42773] = 16'hb89b;
mem_array[42772] = 16'h3e9b;
mem_array[42775] = 16'h14e1;
mem_array[42774] = 16'h3b2d;
mem_array[42777] = 16'h7eb1;
mem_array[42776] = 16'hbed4;
mem_array[42779] = 16'h0221;
mem_array[42778] = 16'hbfc8;
mem_array[42781] = 16'h8bc9;
mem_array[42780] = 16'h3dc4;
mem_array[42783] = 16'h721d;
mem_array[42782] = 16'h3c40;
mem_array[42785] = 16'h3535;
mem_array[42784] = 16'hbdb1;
mem_array[42787] = 16'h862b;
mem_array[42786] = 16'hbfac;
mem_array[42789] = 16'hacce;
mem_array[42788] = 16'hbf56;
mem_array[42791] = 16'hb002;
mem_array[42790] = 16'hbeb4;
mem_array[42793] = 16'h630a;
mem_array[42792] = 16'h3f06;
mem_array[42795] = 16'h5307;
mem_array[42794] = 16'hbe1c;
mem_array[42797] = 16'hd2a1;
mem_array[42796] = 16'hbe8c;
mem_array[42799] = 16'h0147;
mem_array[42798] = 16'hbf5e;
mem_array[42801] = 16'he954;
mem_array[42800] = 16'h3d7e;
mem_array[42803] = 16'h560c;
mem_array[42802] = 16'h3cca;
mem_array[42805] = 16'h0b8c;
mem_array[42804] = 16'hc001;
mem_array[42807] = 16'hbf3c;
mem_array[42806] = 16'hbf72;
mem_array[42809] = 16'h72a1;
mem_array[42808] = 16'h3eae;
mem_array[42811] = 16'hc4c4;
mem_array[42810] = 16'hbd01;
mem_array[42813] = 16'h5bcc;
mem_array[42812] = 16'hbee4;
mem_array[42815] = 16'h209f;
mem_array[42814] = 16'hbed8;
mem_array[42817] = 16'h715c;
mem_array[42816] = 16'h3d2c;
mem_array[42819] = 16'h4b4d;
mem_array[42818] = 16'hbe63;
mem_array[42821] = 16'h29e5;
mem_array[42820] = 16'hbd98;
mem_array[42823] = 16'ha50e;
mem_array[42822] = 16'h3e8c;
mem_array[42825] = 16'h7b5f;
mem_array[42824] = 16'hbf09;
mem_array[42827] = 16'h43c8;
mem_array[42826] = 16'hbe8e;
mem_array[42829] = 16'h531a;
mem_array[42828] = 16'hbe26;
mem_array[42831] = 16'ha1fd;
mem_array[42830] = 16'h3d6d;
mem_array[42833] = 16'h6b97;
mem_array[42832] = 16'h3ede;
mem_array[42835] = 16'hcf16;
mem_array[42834] = 16'h3d95;
mem_array[42837] = 16'he47c;
mem_array[42836] = 16'hbf1d;
mem_array[42839] = 16'h63d7;
mem_array[42838] = 16'hbeff;
mem_array[42841] = 16'h2d76;
mem_array[42840] = 16'h3eb3;
mem_array[42843] = 16'he50d;
mem_array[42842] = 16'h3eca;
mem_array[42845] = 16'ha70c;
mem_array[42844] = 16'h3e65;
mem_array[42847] = 16'h1999;
mem_array[42846] = 16'hbfc2;
mem_array[42849] = 16'hfd8e;
mem_array[42848] = 16'hbfd6;
mem_array[42851] = 16'h37e9;
mem_array[42850] = 16'hbea0;
mem_array[42853] = 16'h86df;
mem_array[42852] = 16'h3e91;
mem_array[42855] = 16'hee6f;
mem_array[42854] = 16'h3e8b;
mem_array[42857] = 16'h428f;
mem_array[42856] = 16'h3c5b;
mem_array[42859] = 16'h13a4;
mem_array[42858] = 16'h3e90;
mem_array[42861] = 16'h5b12;
mem_array[42860] = 16'h3d8b;
mem_array[42863] = 16'he76c;
mem_array[42862] = 16'hbd75;
mem_array[42865] = 16'h588b;
mem_array[42864] = 16'hbfeb;
mem_array[42867] = 16'he5c9;
mem_array[42866] = 16'hbf84;
mem_array[42869] = 16'h7658;
mem_array[42868] = 16'h3e66;
mem_array[42871] = 16'h7b5c;
mem_array[42870] = 16'h3d04;
mem_array[42873] = 16'heb86;
mem_array[42872] = 16'h3e18;
mem_array[42875] = 16'h7073;
mem_array[42874] = 16'hbe13;
mem_array[42877] = 16'hca80;
mem_array[42876] = 16'h3dd3;
mem_array[42879] = 16'ha187;
mem_array[42878] = 16'hbeb4;
mem_array[42881] = 16'h7330;
mem_array[42880] = 16'hbd4f;
mem_array[42883] = 16'h9241;
mem_array[42882] = 16'hbc0a;
mem_array[42885] = 16'h7791;
mem_array[42884] = 16'hbf33;
mem_array[42887] = 16'h53f6;
mem_array[42886] = 16'hbe18;
mem_array[42889] = 16'h5cc8;
mem_array[42888] = 16'hbec8;
mem_array[42891] = 16'h1d0a;
mem_array[42890] = 16'h3df6;
mem_array[42893] = 16'h9fec;
mem_array[42892] = 16'h3e43;
mem_array[42895] = 16'h9a56;
mem_array[42894] = 16'h3d92;
mem_array[42897] = 16'hc38c;
mem_array[42896] = 16'hbe90;
mem_array[42899] = 16'hbeaa;
mem_array[42898] = 16'hbf53;
mem_array[42901] = 16'h585b;
mem_array[42900] = 16'h3c2a;
mem_array[42903] = 16'h776a;
mem_array[42902] = 16'hbe1a;
mem_array[42905] = 16'h8945;
mem_array[42904] = 16'h3ed5;
mem_array[42907] = 16'he037;
mem_array[42906] = 16'hbf75;
mem_array[42909] = 16'hf36d;
mem_array[42908] = 16'hbff9;
mem_array[42911] = 16'h2108;
mem_array[42910] = 16'hbde8;
mem_array[42913] = 16'h2c89;
mem_array[42912] = 16'hbea9;
mem_array[42915] = 16'h0e81;
mem_array[42914] = 16'h3eaa;
mem_array[42917] = 16'h7081;
mem_array[42916] = 16'hbdb2;
mem_array[42919] = 16'h602a;
mem_array[42918] = 16'hbf72;
mem_array[42921] = 16'h8511;
mem_array[42920] = 16'h3d55;
mem_array[42923] = 16'hd09c;
mem_array[42922] = 16'h3cae;
mem_array[42925] = 16'h7c46;
mem_array[42924] = 16'hbfc6;
mem_array[42927] = 16'h0ab9;
mem_array[42926] = 16'hbffe;
mem_array[42929] = 16'h8235;
mem_array[42928] = 16'hbf39;
mem_array[42931] = 16'h690d;
mem_array[42930] = 16'hbe9e;
mem_array[42933] = 16'h9b92;
mem_array[42932] = 16'h3f36;
mem_array[42935] = 16'ha4f7;
mem_array[42934] = 16'hbe00;
mem_array[42937] = 16'h4c91;
mem_array[42936] = 16'hbd43;
mem_array[42939] = 16'h66c6;
mem_array[42938] = 16'h3e7d;
mem_array[42941] = 16'ha323;
mem_array[42940] = 16'h3c9c;
mem_array[42943] = 16'h26f4;
mem_array[42942] = 16'h3e5f;
mem_array[42945] = 16'hd5c6;
mem_array[42944] = 16'hbe88;
mem_array[42947] = 16'h5da7;
mem_array[42946] = 16'h3ef6;
mem_array[42949] = 16'hdb5b;
mem_array[42948] = 16'hbea0;
mem_array[42951] = 16'hd67d;
mem_array[42950] = 16'h3e97;
mem_array[42953] = 16'h5cc3;
mem_array[42952] = 16'h3edc;
mem_array[42955] = 16'h6e6b;
mem_array[42954] = 16'hbd54;
mem_array[42957] = 16'hf68e;
mem_array[42956] = 16'h3eb4;
mem_array[42959] = 16'hd4fd;
mem_array[42958] = 16'hbf31;
mem_array[42961] = 16'h1d8e;
mem_array[42960] = 16'hbf6a;
mem_array[42963] = 16'h18ea;
mem_array[42962] = 16'h3e9d;
mem_array[42965] = 16'h6445;
mem_array[42964] = 16'h3e84;
mem_array[42967] = 16'he397;
mem_array[42966] = 16'hc023;
mem_array[42969] = 16'h43e0;
mem_array[42968] = 16'hbfd0;
mem_array[42971] = 16'hddc8;
mem_array[42970] = 16'hbf07;
mem_array[42973] = 16'h368a;
mem_array[42972] = 16'h3e87;
mem_array[42975] = 16'h2743;
mem_array[42974] = 16'h3cd1;
mem_array[42977] = 16'h594f;
mem_array[42976] = 16'h3e94;
mem_array[42979] = 16'h0055;
mem_array[42978] = 16'hbfdb;
mem_array[42981] = 16'hc3f2;
mem_array[42980] = 16'hbcfe;
mem_array[42983] = 16'h5260;
mem_array[42982] = 16'hbda7;
mem_array[42985] = 16'h7711;
mem_array[42984] = 16'hbfa0;
mem_array[42987] = 16'hb591;
mem_array[42986] = 16'hbf67;
mem_array[42989] = 16'h17bd;
mem_array[42988] = 16'h3e30;
mem_array[42991] = 16'hf59b;
mem_array[42990] = 16'hbe2d;
mem_array[42993] = 16'h21b6;
mem_array[42992] = 16'hbf08;
mem_array[42995] = 16'h021d;
mem_array[42994] = 16'hbee3;
mem_array[42997] = 16'hbcc7;
mem_array[42996] = 16'h3bbc;
mem_array[42999] = 16'h037a;
mem_array[42998] = 16'hbe8c;
mem_array[43001] = 16'h9534;
mem_array[43000] = 16'hbef6;
mem_array[43003] = 16'h77a3;
mem_array[43002] = 16'h3ea7;
mem_array[43005] = 16'h7278;
mem_array[43004] = 16'hbf51;
mem_array[43007] = 16'h057c;
mem_array[43006] = 16'h3e99;
mem_array[43009] = 16'h23eb;
mem_array[43008] = 16'hbe1d;
mem_array[43011] = 16'h66bb;
mem_array[43010] = 16'h3ee0;
mem_array[43013] = 16'h0411;
mem_array[43012] = 16'h3eca;
mem_array[43015] = 16'h56fe;
mem_array[43014] = 16'hbe80;
mem_array[43017] = 16'h5aed;
mem_array[43016] = 16'h3e7a;
mem_array[43019] = 16'hfac6;
mem_array[43018] = 16'hbf9e;
mem_array[43021] = 16'h9039;
mem_array[43020] = 16'hbf1d;
mem_array[43023] = 16'h42d0;
mem_array[43022] = 16'h3e8b;
mem_array[43025] = 16'hf522;
mem_array[43024] = 16'hbe2e;
mem_array[43027] = 16'hd317;
mem_array[43026] = 16'hc030;
mem_array[43029] = 16'haa3e;
mem_array[43028] = 16'hbed4;
mem_array[43031] = 16'h41eb;
mem_array[43030] = 16'hbeb9;
mem_array[43033] = 16'h0c43;
mem_array[43032] = 16'h3e57;
mem_array[43035] = 16'h92cd;
mem_array[43034] = 16'h3dd2;
mem_array[43037] = 16'h721b;
mem_array[43036] = 16'h3e14;
mem_array[43039] = 16'hb624;
mem_array[43038] = 16'hbf83;
mem_array[43041] = 16'h6600;
mem_array[43040] = 16'hba0b;
mem_array[43043] = 16'hee81;
mem_array[43042] = 16'hbd2b;
mem_array[43045] = 16'h71ba;
mem_array[43044] = 16'hc013;
mem_array[43047] = 16'h2f21;
mem_array[43046] = 16'hbebf;
mem_array[43049] = 16'ha3ff;
mem_array[43048] = 16'hbe9f;
mem_array[43051] = 16'h1356;
mem_array[43050] = 16'hba50;
mem_array[43053] = 16'h3f89;
mem_array[43052] = 16'hbf1c;
mem_array[43055] = 16'h2d00;
mem_array[43054] = 16'h3e8b;
mem_array[43057] = 16'h6ca5;
mem_array[43056] = 16'hbe5c;
mem_array[43059] = 16'hb6f4;
mem_array[43058] = 16'hbea4;
mem_array[43061] = 16'h8aee;
mem_array[43060] = 16'hbebe;
mem_array[43063] = 16'h675a;
mem_array[43062] = 16'h3f63;
mem_array[43065] = 16'hbe49;
mem_array[43064] = 16'hbdec;
mem_array[43067] = 16'h451a;
mem_array[43066] = 16'h3d88;
mem_array[43069] = 16'h5dcb;
mem_array[43068] = 16'hbe8f;
mem_array[43071] = 16'hbebb;
mem_array[43070] = 16'h3bbc;
mem_array[43073] = 16'hf759;
mem_array[43072] = 16'h3e8d;
mem_array[43075] = 16'h5685;
mem_array[43074] = 16'h3f3d;
mem_array[43077] = 16'h7284;
mem_array[43076] = 16'h3f12;
mem_array[43079] = 16'hb247;
mem_array[43078] = 16'hbf7e;
mem_array[43081] = 16'h6c91;
mem_array[43080] = 16'hbf35;
mem_array[43083] = 16'hca12;
mem_array[43082] = 16'hbe8a;
mem_array[43085] = 16'h0498;
mem_array[43084] = 16'hbee1;
mem_array[43087] = 16'h9ad2;
mem_array[43086] = 16'hc029;
mem_array[43089] = 16'h211a;
mem_array[43088] = 16'h3e19;
mem_array[43091] = 16'hc04a;
mem_array[43090] = 16'hbf6a;
mem_array[43093] = 16'hba6d;
mem_array[43092] = 16'h3eb2;
mem_array[43095] = 16'h3a3e;
mem_array[43094] = 16'h3e6a;
mem_array[43097] = 16'h979a;
mem_array[43096] = 16'hbed1;
mem_array[43099] = 16'he646;
mem_array[43098] = 16'hbf44;
mem_array[43101] = 16'h18d1;
mem_array[43100] = 16'h3b19;
mem_array[43103] = 16'hfeb0;
mem_array[43102] = 16'h3d8f;
mem_array[43105] = 16'hf40f;
mem_array[43104] = 16'hbffd;
mem_array[43107] = 16'h5913;
mem_array[43106] = 16'h3ec3;
mem_array[43109] = 16'h55cf;
mem_array[43108] = 16'hbe67;
mem_array[43111] = 16'he0c4;
mem_array[43110] = 16'h3ea2;
mem_array[43113] = 16'h6787;
mem_array[43112] = 16'hbf01;
mem_array[43115] = 16'h0e71;
mem_array[43114] = 16'h3e65;
mem_array[43117] = 16'hf771;
mem_array[43116] = 16'h3e50;
mem_array[43119] = 16'h3a1a;
mem_array[43118] = 16'hbf30;
mem_array[43121] = 16'h0dc3;
mem_array[43120] = 16'hbd6e;
mem_array[43123] = 16'hc0e6;
mem_array[43122] = 16'h3e95;
mem_array[43125] = 16'he8c7;
mem_array[43124] = 16'hbd07;
mem_array[43127] = 16'h183d;
mem_array[43126] = 16'hbdf9;
mem_array[43129] = 16'h06d0;
mem_array[43128] = 16'h3dc9;
mem_array[43131] = 16'h1bde;
mem_array[43130] = 16'h3e97;
mem_array[43133] = 16'h6fc2;
mem_array[43132] = 16'h3e01;
mem_array[43135] = 16'h445b;
mem_array[43134] = 16'h3f1f;
mem_array[43137] = 16'h2d82;
mem_array[43136] = 16'h3f0e;
mem_array[43139] = 16'h9437;
mem_array[43138] = 16'hbee2;
mem_array[43141] = 16'h7848;
mem_array[43140] = 16'hbeec;
mem_array[43143] = 16'h95aa;
mem_array[43142] = 16'h3f22;
mem_array[43145] = 16'haca6;
mem_array[43144] = 16'hbe88;
mem_array[43147] = 16'h1878;
mem_array[43146] = 16'hc02d;
mem_array[43149] = 16'haa46;
mem_array[43148] = 16'hbec0;
mem_array[43151] = 16'hd8e5;
mem_array[43150] = 16'hbf3a;
mem_array[43153] = 16'hce64;
mem_array[43152] = 16'h4008;
mem_array[43155] = 16'hefad;
mem_array[43154] = 16'h3ef6;
mem_array[43157] = 16'hc25d;
mem_array[43156] = 16'hbe52;
mem_array[43159] = 16'h56c0;
mem_array[43158] = 16'hbee6;
mem_array[43161] = 16'ha888;
mem_array[43160] = 16'h3c97;
mem_array[43163] = 16'h60ea;
mem_array[43162] = 16'hbc0e;
mem_array[43165] = 16'ha502;
mem_array[43164] = 16'hbfef;
mem_array[43167] = 16'h945c;
mem_array[43166] = 16'hbec0;
mem_array[43169] = 16'h214d;
mem_array[43168] = 16'hbe67;
mem_array[43171] = 16'h42a5;
mem_array[43170] = 16'hbecf;
mem_array[43173] = 16'h0144;
mem_array[43172] = 16'hbeef;
mem_array[43175] = 16'h1ca7;
mem_array[43174] = 16'hbedc;
mem_array[43177] = 16'h18b4;
mem_array[43176] = 16'hbe9d;
mem_array[43179] = 16'ha153;
mem_array[43178] = 16'hbec7;
mem_array[43181] = 16'hb76c;
mem_array[43180] = 16'hbf0a;
mem_array[43183] = 16'h9df9;
mem_array[43182] = 16'h3e6f;
mem_array[43185] = 16'hbf3b;
mem_array[43184] = 16'hbf55;
mem_array[43187] = 16'h2416;
mem_array[43186] = 16'h3eb6;
mem_array[43189] = 16'h5fff;
mem_array[43188] = 16'h3e83;
mem_array[43191] = 16'ha5a0;
mem_array[43190] = 16'hbea8;
mem_array[43193] = 16'h7fda;
mem_array[43192] = 16'h3f43;
mem_array[43195] = 16'h9b96;
mem_array[43194] = 16'h3ebd;
mem_array[43197] = 16'hdcab;
mem_array[43196] = 16'hbe01;
mem_array[43199] = 16'h44d5;
mem_array[43198] = 16'hbfd5;
mem_array[43201] = 16'h7546;
mem_array[43200] = 16'hbe1c;
mem_array[43203] = 16'h4df7;
mem_array[43202] = 16'h3eba;
mem_array[43205] = 16'h502e;
mem_array[43204] = 16'hbe9b;
mem_array[43207] = 16'h86bc;
mem_array[43206] = 16'hbfb8;
mem_array[43209] = 16'h0a00;
mem_array[43208] = 16'h3eb8;
mem_array[43211] = 16'h56ee;
mem_array[43210] = 16'h3e42;
mem_array[43213] = 16'h08dc;
mem_array[43212] = 16'h3e1a;
mem_array[43215] = 16'h4716;
mem_array[43214] = 16'h3f37;
mem_array[43217] = 16'hb5d9;
mem_array[43216] = 16'hbe17;
mem_array[43219] = 16'h5c5e;
mem_array[43218] = 16'hbed6;
mem_array[43221] = 16'h0cd2;
mem_array[43220] = 16'hbca5;
mem_array[43223] = 16'hb9e8;
mem_array[43222] = 16'hbb89;
mem_array[43225] = 16'hf2b6;
mem_array[43224] = 16'hbf9f;
mem_array[43227] = 16'hc6f1;
mem_array[43226] = 16'hbf84;
mem_array[43229] = 16'h972a;
mem_array[43228] = 16'h3ed3;
mem_array[43231] = 16'hd4e5;
mem_array[43230] = 16'hbe09;
mem_array[43233] = 16'hb3e3;
mem_array[43232] = 16'h3f48;
mem_array[43235] = 16'h0e39;
mem_array[43234] = 16'hbeed;
mem_array[43237] = 16'h3177;
mem_array[43236] = 16'h3c29;
mem_array[43239] = 16'h737d;
mem_array[43238] = 16'hbf20;
mem_array[43241] = 16'h976d;
mem_array[43240] = 16'h3edf;
mem_array[43243] = 16'h1091;
mem_array[43242] = 16'hbe08;
mem_array[43245] = 16'hcca9;
mem_array[43244] = 16'hbdf7;
mem_array[43247] = 16'hf074;
mem_array[43246] = 16'h3eb6;
mem_array[43249] = 16'h7ce4;
mem_array[43248] = 16'h3ea5;
mem_array[43251] = 16'hee24;
mem_array[43250] = 16'hbf85;
mem_array[43253] = 16'he944;
mem_array[43252] = 16'h3d1f;
mem_array[43255] = 16'h4d07;
mem_array[43254] = 16'hbe52;
mem_array[43257] = 16'h34ea;
mem_array[43256] = 16'hbe78;
mem_array[43259] = 16'h02c7;
mem_array[43258] = 16'hbfb6;
mem_array[43261] = 16'h108e;
mem_array[43260] = 16'hbe41;
mem_array[43263] = 16'h4742;
mem_array[43262] = 16'h3f40;
mem_array[43265] = 16'h58ad;
mem_array[43264] = 16'hbee6;
mem_array[43267] = 16'h8380;
mem_array[43266] = 16'hbf65;
mem_array[43269] = 16'h9945;
mem_array[43268] = 16'hbe49;
mem_array[43271] = 16'hb401;
mem_array[43270] = 16'hbdd4;
mem_array[43273] = 16'h8be4;
mem_array[43272] = 16'hbedb;
mem_array[43275] = 16'h3078;
mem_array[43274] = 16'h3f21;
mem_array[43277] = 16'h6f9d;
mem_array[43276] = 16'hbebc;
mem_array[43279] = 16'h08ec;
mem_array[43278] = 16'h3d9d;
mem_array[43281] = 16'hc644;
mem_array[43280] = 16'hbcf2;
mem_array[43283] = 16'h9a44;
mem_array[43282] = 16'hbdb5;
mem_array[43285] = 16'he6de;
mem_array[43284] = 16'hbfc0;
mem_array[43287] = 16'h2220;
mem_array[43286] = 16'hbf84;
mem_array[43289] = 16'hf31d;
mem_array[43288] = 16'hbd6a;
mem_array[43291] = 16'h4e77;
mem_array[43290] = 16'hbf08;
mem_array[43293] = 16'hd2a7;
mem_array[43292] = 16'hbe86;
mem_array[43295] = 16'h3d79;
mem_array[43294] = 16'hbf24;
mem_array[43297] = 16'hbb7b;
mem_array[43296] = 16'hbea2;
mem_array[43299] = 16'h9084;
mem_array[43298] = 16'hbef5;
mem_array[43301] = 16'h216c;
mem_array[43300] = 16'h3df1;
mem_array[43303] = 16'h4fee;
mem_array[43302] = 16'h3ee1;
mem_array[43305] = 16'h0b5c;
mem_array[43304] = 16'hbcd1;
mem_array[43307] = 16'h885a;
mem_array[43306] = 16'h3f06;
mem_array[43309] = 16'hfc14;
mem_array[43308] = 16'hbf0f;
mem_array[43311] = 16'h7612;
mem_array[43310] = 16'hbf94;
mem_array[43313] = 16'ha11d;
mem_array[43312] = 16'h3d1b;
mem_array[43315] = 16'h556f;
mem_array[43314] = 16'h3e98;
mem_array[43317] = 16'h00af;
mem_array[43316] = 16'hbee1;
mem_array[43319] = 16'h6d22;
mem_array[43318] = 16'hbfcc;
mem_array[43321] = 16'h0d1e;
mem_array[43320] = 16'h3ecf;
mem_array[43323] = 16'hc70f;
mem_array[43322] = 16'h3dab;
mem_array[43325] = 16'hf7b1;
mem_array[43324] = 16'hbfa0;
mem_array[43327] = 16'h6849;
mem_array[43326] = 16'hbf7b;
mem_array[43329] = 16'h8c48;
mem_array[43328] = 16'h3d5b;
mem_array[43331] = 16'h38bf;
mem_array[43330] = 16'hbe21;
mem_array[43333] = 16'hec49;
mem_array[43332] = 16'hbf1f;
mem_array[43335] = 16'hfa23;
mem_array[43334] = 16'h3f22;
mem_array[43337] = 16'hba15;
mem_array[43336] = 16'hbee9;
mem_array[43339] = 16'h339a;
mem_array[43338] = 16'h3e27;
mem_array[43341] = 16'hb3fa;
mem_array[43340] = 16'hbd0e;
mem_array[43343] = 16'h1cf4;
mem_array[43342] = 16'h3a86;
mem_array[43345] = 16'h2165;
mem_array[43344] = 16'hbf56;
mem_array[43347] = 16'h8d17;
mem_array[43346] = 16'hbf26;
mem_array[43349] = 16'hcf40;
mem_array[43348] = 16'hbd9f;
mem_array[43351] = 16'hbd28;
mem_array[43350] = 16'hbf8a;
mem_array[43353] = 16'h014d;
mem_array[43352] = 16'hbe1a;
mem_array[43355] = 16'hdebf;
mem_array[43354] = 16'hbe6b;
mem_array[43357] = 16'h019d;
mem_array[43356] = 16'hbf8a;
mem_array[43359] = 16'h9fa5;
mem_array[43358] = 16'hbf81;
mem_array[43361] = 16'h5931;
mem_array[43360] = 16'h3ec0;
mem_array[43363] = 16'h2bf3;
mem_array[43362] = 16'h3f7e;
mem_array[43365] = 16'h2556;
mem_array[43364] = 16'hbd64;
mem_array[43367] = 16'h02c7;
mem_array[43366] = 16'h3f39;
mem_array[43369] = 16'h06e2;
mem_array[43368] = 16'hbf6d;
mem_array[43371] = 16'hb481;
mem_array[43370] = 16'hbf30;
mem_array[43373] = 16'hf09d;
mem_array[43372] = 16'h3e2b;
mem_array[43375] = 16'hb310;
mem_array[43374] = 16'h3ef1;
mem_array[43377] = 16'hc09a;
mem_array[43376] = 16'hbe5b;
mem_array[43379] = 16'hda1c;
mem_array[43378] = 16'hbefc;
mem_array[43381] = 16'h8f12;
mem_array[43380] = 16'hbf98;
mem_array[43383] = 16'hcba3;
mem_array[43382] = 16'hbebd;
mem_array[43385] = 16'h247f;
mem_array[43384] = 16'hbf8b;
mem_array[43387] = 16'he506;
mem_array[43386] = 16'hbf9d;
mem_array[43389] = 16'h0281;
mem_array[43388] = 16'h3ceb;
mem_array[43391] = 16'h43aa;
mem_array[43390] = 16'hbf0b;
mem_array[43393] = 16'hf608;
mem_array[43392] = 16'hbf87;
mem_array[43395] = 16'ha9a2;
mem_array[43394] = 16'hbf91;
mem_array[43397] = 16'hdf6c;
mem_array[43396] = 16'hbe71;
mem_array[43399] = 16'h7e7b;
mem_array[43398] = 16'hbd80;
mem_array[43401] = 16'he63b;
mem_array[43400] = 16'hbd3d;
mem_array[43403] = 16'hd4c5;
mem_array[43402] = 16'h3b73;
mem_array[43405] = 16'h4464;
mem_array[43404] = 16'h3f01;
mem_array[43407] = 16'h3eb8;
mem_array[43406] = 16'hbe05;
mem_array[43409] = 16'hd77d;
mem_array[43408] = 16'h3e71;
mem_array[43411] = 16'h9a74;
mem_array[43410] = 16'hbf8b;
mem_array[43413] = 16'h3c69;
mem_array[43412] = 16'hbe46;
mem_array[43415] = 16'h94f9;
mem_array[43414] = 16'h3eca;
mem_array[43417] = 16'hc428;
mem_array[43416] = 16'hbe2a;
mem_array[43419] = 16'he758;
mem_array[43418] = 16'hbe8e;
mem_array[43421] = 16'h663b;
mem_array[43420] = 16'h3f8f;
mem_array[43423] = 16'h9b97;
mem_array[43422] = 16'h3f14;
mem_array[43425] = 16'h7dd6;
mem_array[43424] = 16'hbd64;
mem_array[43427] = 16'hacb6;
mem_array[43426] = 16'h3db5;
mem_array[43429] = 16'hfc02;
mem_array[43428] = 16'h3e94;
mem_array[43431] = 16'haaf2;
mem_array[43430] = 16'hbea8;
mem_array[43433] = 16'h5634;
mem_array[43432] = 16'hbf81;
mem_array[43435] = 16'h2da8;
mem_array[43434] = 16'hbd97;
mem_array[43437] = 16'hb4f4;
mem_array[43436] = 16'hbd9f;
mem_array[43439] = 16'h5825;
mem_array[43438] = 16'h3e4e;
mem_array[43441] = 16'h8b16;
mem_array[43440] = 16'hbdb3;
mem_array[43443] = 16'h31ab;
mem_array[43442] = 16'h3d30;
mem_array[43445] = 16'h5380;
mem_array[43444] = 16'hbf09;
mem_array[43447] = 16'hf227;
mem_array[43446] = 16'hbec0;
mem_array[43449] = 16'h5730;
mem_array[43448] = 16'hbebb;
mem_array[43451] = 16'h6e81;
mem_array[43450] = 16'hbcd4;
mem_array[43453] = 16'hfe8f;
mem_array[43452] = 16'hbc33;
mem_array[43455] = 16'he7cf;
mem_array[43454] = 16'h3d07;
mem_array[43457] = 16'h9905;
mem_array[43456] = 16'h3d7a;
mem_array[43459] = 16'hcdac;
mem_array[43458] = 16'hbddb;
mem_array[43461] = 16'h9a48;
mem_array[43460] = 16'hbd27;
mem_array[43463] = 16'hcbcd;
mem_array[43462] = 16'hbd34;
mem_array[43465] = 16'ha0a7;
mem_array[43464] = 16'h3e12;
mem_array[43467] = 16'h869a;
mem_array[43466] = 16'h3f3b;
mem_array[43469] = 16'h2694;
mem_array[43468] = 16'h3f05;
mem_array[43471] = 16'h9b81;
mem_array[43470] = 16'hbfc6;
mem_array[43473] = 16'h42d3;
mem_array[43472] = 16'hbc65;
mem_array[43475] = 16'hdf78;
mem_array[43474] = 16'hbe8d;
mem_array[43477] = 16'hc108;
mem_array[43476] = 16'hbef1;
mem_array[43479] = 16'h89e0;
mem_array[43478] = 16'hbf3b;
mem_array[43481] = 16'hb116;
mem_array[43480] = 16'hbe9a;
mem_array[43483] = 16'ha837;
mem_array[43482] = 16'h3fbc;
mem_array[43485] = 16'h6799;
mem_array[43484] = 16'h3c82;
mem_array[43487] = 16'h3be4;
mem_array[43486] = 16'hbe3d;
mem_array[43489] = 16'h1d5f;
mem_array[43488] = 16'h3ed0;
mem_array[43491] = 16'he7a7;
mem_array[43490] = 16'h3ee4;
mem_array[43493] = 16'h1205;
mem_array[43492] = 16'h3eaf;
mem_array[43495] = 16'h56d1;
mem_array[43494] = 16'hbe20;
mem_array[43497] = 16'hf515;
mem_array[43496] = 16'hbd7a;
mem_array[43499] = 16'h6748;
mem_array[43498] = 16'hbf3a;
mem_array[43501] = 16'h4714;
mem_array[43500] = 16'hbd15;
mem_array[43503] = 16'h4c02;
mem_array[43502] = 16'hbc94;
mem_array[43505] = 16'hd049;
mem_array[43504] = 16'h3e9e;
mem_array[43507] = 16'ha709;
mem_array[43506] = 16'hbd9c;
mem_array[43509] = 16'h1057;
mem_array[43508] = 16'hbb7e;
mem_array[43511] = 16'h8c43;
mem_array[43510] = 16'hbd61;
mem_array[43513] = 16'hd2a7;
mem_array[43512] = 16'hbdb0;
mem_array[43515] = 16'he21e;
mem_array[43514] = 16'h3d53;
mem_array[43517] = 16'hd87e;
mem_array[43516] = 16'h3dc0;
mem_array[43519] = 16'hab10;
mem_array[43518] = 16'hbd32;
mem_array[43521] = 16'h563e;
mem_array[43520] = 16'hbd22;
mem_array[43523] = 16'ha0f1;
mem_array[43522] = 16'hbd87;
mem_array[43525] = 16'h31a9;
mem_array[43524] = 16'hbd59;
mem_array[43527] = 16'h5635;
mem_array[43526] = 16'h3f48;
mem_array[43529] = 16'h1ee1;
mem_array[43528] = 16'h3ef4;
mem_array[43531] = 16'h4d1a;
mem_array[43530] = 16'h3e32;
mem_array[43533] = 16'h3770;
mem_array[43532] = 16'hbc89;
mem_array[43535] = 16'h77aa;
mem_array[43534] = 16'hbdc3;
mem_array[43537] = 16'h8107;
mem_array[43536] = 16'h3f09;
mem_array[43539] = 16'ha2b9;
mem_array[43538] = 16'hbdc5;
mem_array[43541] = 16'h699a;
mem_array[43540] = 16'hbd99;
mem_array[43543] = 16'haf5c;
mem_array[43542] = 16'hbf5c;
mem_array[43545] = 16'h86bb;
mem_array[43544] = 16'hbcb9;
mem_array[43547] = 16'h1876;
mem_array[43546] = 16'hbea0;
mem_array[43549] = 16'hc359;
mem_array[43548] = 16'h3f0b;
mem_array[43551] = 16'hee6e;
mem_array[43550] = 16'hbdb8;
mem_array[43553] = 16'hd889;
mem_array[43552] = 16'hbe32;
mem_array[43555] = 16'hd9dd;
mem_array[43554] = 16'hbd6f;
mem_array[43557] = 16'hdf76;
mem_array[43556] = 16'h3ada;
mem_array[43559] = 16'h15f2;
mem_array[43558] = 16'hbd90;
mem_array[43561] = 16'h1baa;
mem_array[43560] = 16'h3d2a;
mem_array[43563] = 16'h0d71;
mem_array[43562] = 16'h3de4;
mem_array[43565] = 16'h923e;
mem_array[43564] = 16'h3f3d;
mem_array[43567] = 16'h6a3d;
mem_array[43566] = 16'h3d8c;
mem_array[43569] = 16'h6783;
mem_array[43568] = 16'h3ce5;
mem_array[43571] = 16'h0282;
mem_array[43570] = 16'h39dc;
mem_array[43573] = 16'h859b;
mem_array[43572] = 16'h3d9e;
mem_array[43575] = 16'h0b8b;
mem_array[43574] = 16'hbc87;
mem_array[43577] = 16'h8b7a;
mem_array[43576] = 16'h3da1;
mem_array[43579] = 16'h5769;
mem_array[43578] = 16'hbd50;
mem_array[43581] = 16'h4388;
mem_array[43580] = 16'h3d0c;
mem_array[43583] = 16'h0c1c;
mem_array[43582] = 16'h3d7f;
mem_array[43585] = 16'h53e1;
mem_array[43584] = 16'h3d2d;
mem_array[43587] = 16'h7457;
mem_array[43586] = 16'h3f5c;
mem_array[43589] = 16'hc154;
mem_array[43588] = 16'h3f1c;
mem_array[43591] = 16'hc4cb;
mem_array[43590] = 16'h3e85;
mem_array[43593] = 16'h5560;
mem_array[43592] = 16'h3d83;
mem_array[43595] = 16'h4f0c;
mem_array[43594] = 16'h3c94;
mem_array[43597] = 16'h7c88;
mem_array[43596] = 16'hbeaf;
mem_array[43599] = 16'h23a9;
mem_array[43598] = 16'h3b83;
mem_array[43601] = 16'h75bb;
mem_array[43600] = 16'hbd7a;
mem_array[43603] = 16'hd04b;
mem_array[43602] = 16'hbe89;
mem_array[43605] = 16'haa9a;
mem_array[43604] = 16'h3c51;
mem_array[43607] = 16'hc76d;
mem_array[43606] = 16'hbf50;
mem_array[43609] = 16'hc41d;
mem_array[43608] = 16'h3f42;
mem_array[43611] = 16'hc586;
mem_array[43610] = 16'h3d8a;
mem_array[43613] = 16'h5719;
mem_array[43612] = 16'h3f2f;
mem_array[43615] = 16'h865e;
mem_array[43614] = 16'h3d5f;
mem_array[43617] = 16'ha8e3;
mem_array[43616] = 16'hbd73;
mem_array[43619] = 16'h966b;
mem_array[43618] = 16'hbdb8;
mem_array[43621] = 16'hae7a;
mem_array[43620] = 16'hbd81;
mem_array[43623] = 16'h8d49;
mem_array[43622] = 16'hbd88;
mem_array[43625] = 16'hdbbc;
mem_array[43624] = 16'h3dbf;
mem_array[43627] = 16'h6db0;
mem_array[43626] = 16'h3d26;
mem_array[43629] = 16'hfe22;
mem_array[43628] = 16'hbca0;
mem_array[43631] = 16'h62ae;
mem_array[43630] = 16'hbaa4;
mem_array[43633] = 16'h87b6;
mem_array[43632] = 16'hbd2d;
mem_array[43635] = 16'hc34a;
mem_array[43634] = 16'hbc06;
mem_array[43637] = 16'h684f;
mem_array[43636] = 16'h3d8f;
mem_array[43639] = 16'hcca3;
mem_array[43638] = 16'hbcd8;
mem_array[43641] = 16'hb97d;
mem_array[43640] = 16'hba6d;
mem_array[43643] = 16'hf4ea;
mem_array[43642] = 16'hbd13;
mem_array[43645] = 16'h5046;
mem_array[43644] = 16'h3bb7;
mem_array[43647] = 16'h4af6;
mem_array[43646] = 16'h3db7;
mem_array[43649] = 16'h3854;
mem_array[43648] = 16'hbd3f;
mem_array[43651] = 16'h0fd7;
mem_array[43650] = 16'hbbe8;
mem_array[43653] = 16'hd8e7;
mem_array[43652] = 16'h3d33;
mem_array[43655] = 16'hda88;
mem_array[43654] = 16'h3d74;
mem_array[43657] = 16'h0f5c;
mem_array[43656] = 16'hbd46;
mem_array[43659] = 16'hd226;
mem_array[43658] = 16'hbcb7;
mem_array[43661] = 16'h85f0;
mem_array[43660] = 16'hbb19;
mem_array[43663] = 16'h54bd;
mem_array[43662] = 16'h3d3c;
mem_array[43665] = 16'hf8b0;
mem_array[43664] = 16'hbd98;
mem_array[43667] = 16'h1604;
mem_array[43666] = 16'hbbe0;
mem_array[43669] = 16'ha36e;
mem_array[43668] = 16'h3ca6;
mem_array[43671] = 16'h01fd;
mem_array[43670] = 16'hbd65;
mem_array[43673] = 16'h6b65;
mem_array[43672] = 16'hbde1;
mem_array[43675] = 16'ha478;
mem_array[43674] = 16'h3cbe;
mem_array[43677] = 16'h2000;
mem_array[43676] = 16'h3b88;
mem_array[43679] = 16'h0ac0;
mem_array[43678] = 16'hbd6f;
mem_array[43681] = 16'ha6f9;
mem_array[43680] = 16'hbda1;
mem_array[43683] = 16'h67e2;
mem_array[43682] = 16'h3d67;
mem_array[43685] = 16'hc9db;
mem_array[43684] = 16'h3d9a;
mem_array[43687] = 16'hf644;
mem_array[43686] = 16'hbc1a;
mem_array[43689] = 16'h2d57;
mem_array[43688] = 16'hbdaf;
mem_array[43691] = 16'h6435;
mem_array[43690] = 16'hbdab;
mem_array[43693] = 16'h8eab;
mem_array[43692] = 16'h3d78;
mem_array[43695] = 16'h1100;
mem_array[43694] = 16'h3db6;
mem_array[43697] = 16'h37a1;
mem_array[43696] = 16'hbda3;
mem_array[43699] = 16'h6ae3;
mem_array[43698] = 16'h3d3b;
mem_array[43701] = 16'h02ec;
mem_array[43700] = 16'hbd47;
mem_array[43703] = 16'h7aa9;
mem_array[43702] = 16'h3c24;
mem_array[43705] = 16'h12c0;
mem_array[43704] = 16'hbd22;
mem_array[43707] = 16'h57f6;
mem_array[43706] = 16'h3d47;
mem_array[43709] = 16'hbc1d;
mem_array[43708] = 16'h3d7d;
mem_array[43711] = 16'h44ee;
mem_array[43710] = 16'h3dd5;
mem_array[43713] = 16'h6593;
mem_array[43712] = 16'hbc2d;
mem_array[43715] = 16'h3455;
mem_array[43714] = 16'hbdc4;
mem_array[43717] = 16'h9dd7;
mem_array[43716] = 16'h3ddc;
mem_array[43719] = 16'hca92;
mem_array[43718] = 16'hbd46;
mem_array[43721] = 16'ha6a9;
mem_array[43720] = 16'hbc84;
mem_array[43723] = 16'hddf2;
mem_array[43722] = 16'h3d89;
mem_array[43725] = 16'ha905;
mem_array[43724] = 16'hbd22;
mem_array[43727] = 16'h70ea;
mem_array[43726] = 16'hbcab;
mem_array[43729] = 16'he09f;
mem_array[43728] = 16'hbc05;
mem_array[43731] = 16'hd592;
mem_array[43730] = 16'hbc85;
mem_array[43733] = 16'hbd71;
mem_array[43732] = 16'hbd36;
mem_array[43735] = 16'hd3ba;
mem_array[43734] = 16'h3d82;
mem_array[43737] = 16'h7976;
mem_array[43736] = 16'h3d1b;
mem_array[43739] = 16'h58ac;
mem_array[43738] = 16'h3b0b;
mem_array[43741] = 16'h1c36;
mem_array[43740] = 16'h3c8f;
mem_array[43743] = 16'hd145;
mem_array[43742] = 16'h3c6d;
mem_array[43745] = 16'h8837;
mem_array[43744] = 16'hbd73;
mem_array[43747] = 16'h4c5f;
mem_array[43746] = 16'h3aab;
mem_array[43749] = 16'h4b2b;
mem_array[43748] = 16'h3d75;
mem_array[43751] = 16'hae99;
mem_array[43750] = 16'h3cb9;
mem_array[43753] = 16'h537f;
mem_array[43752] = 16'h3d0d;
mem_array[43755] = 16'h5b7f;
mem_array[43754] = 16'hbc82;
mem_array[43757] = 16'hd327;
mem_array[43756] = 16'hbd18;
mem_array[43759] = 16'h26d3;
mem_array[43758] = 16'h3da6;
mem_array[43761] = 16'h0068;
mem_array[43760] = 16'hbc90;
mem_array[43763] = 16'hb5e6;
mem_array[43762] = 16'h3d0b;
mem_array[43765] = 16'hab52;
mem_array[43764] = 16'h3c63;
mem_array[43767] = 16'hd068;
mem_array[43766] = 16'hbc8e;
mem_array[43769] = 16'hf4a5;
mem_array[43768] = 16'h3cbe;
mem_array[43771] = 16'he513;
mem_array[43770] = 16'h3dba;
mem_array[43773] = 16'h687f;
mem_array[43772] = 16'h3adf;
mem_array[43775] = 16'hdffd;
mem_array[43774] = 16'hbc55;
mem_array[43777] = 16'h3608;
mem_array[43776] = 16'hbc93;
mem_array[43779] = 16'h1563;
mem_array[43778] = 16'h3d90;
mem_array[43781] = 16'h13dd;
mem_array[43780] = 16'hbc70;
mem_array[43783] = 16'hec41;
mem_array[43782] = 16'h3d35;
mem_array[43785] = 16'haa01;
mem_array[43784] = 16'hbd81;
mem_array[43787] = 16'h00bd;
mem_array[43786] = 16'h3d8d;
mem_array[43789] = 16'h5f91;
mem_array[43788] = 16'hbd7a;
mem_array[43791] = 16'h5408;
mem_array[43790] = 16'h3d9b;
mem_array[43793] = 16'hc818;
mem_array[43792] = 16'hbc5a;
mem_array[43795] = 16'hebac;
mem_array[43794] = 16'h3d76;
mem_array[43797] = 16'h95ac;
mem_array[43796] = 16'hbd0c;
mem_array[43799] = 16'h51b2;
mem_array[43798] = 16'hbd43;
mem_array[43801] = 16'h2d96;
mem_array[43800] = 16'h3d30;
mem_array[43803] = 16'h1d3e;
mem_array[43802] = 16'h3d8f;
mem_array[43805] = 16'h035e;
mem_array[43804] = 16'hbcc7;
mem_array[43807] = 16'h322c;
mem_array[43806] = 16'hbcb1;
mem_array[43809] = 16'h69bf;
mem_array[43808] = 16'hbd03;
mem_array[43811] = 16'h3715;
mem_array[43810] = 16'hbcfe;
mem_array[43813] = 16'heec9;
mem_array[43812] = 16'h3de4;
mem_array[43815] = 16'h1e8f;
mem_array[43814] = 16'h3ce7;
mem_array[43817] = 16'h2596;
mem_array[43816] = 16'hbb68;
mem_array[43819] = 16'h355b;
mem_array[43818] = 16'hbd56;
mem_array[43821] = 16'h186f;
mem_array[43820] = 16'h3ce7;
mem_array[43823] = 16'hec8d;
mem_array[43822] = 16'hbc73;
mem_array[43825] = 16'h9f18;
mem_array[43824] = 16'h3d21;
mem_array[43827] = 16'hd5c9;
mem_array[43826] = 16'h3b90;
mem_array[43829] = 16'h65f3;
mem_array[43828] = 16'hbc44;
mem_array[43831] = 16'h1d52;
mem_array[43830] = 16'h3d20;
mem_array[43833] = 16'hed07;
mem_array[43832] = 16'h3d7c;
mem_array[43835] = 16'h1592;
mem_array[43834] = 16'hbc5f;
mem_array[43837] = 16'h666c;
mem_array[43836] = 16'hbd34;
mem_array[43839] = 16'hceb8;
mem_array[43838] = 16'h3d31;
mem_array[43841] = 16'hb19a;
mem_array[43840] = 16'h3d3b;
mem_array[43843] = 16'hf264;
mem_array[43842] = 16'hbdb0;
mem_array[43845] = 16'h3717;
mem_array[43844] = 16'hbd20;
mem_array[43847] = 16'hc3d1;
mem_array[43846] = 16'hbcc8;
mem_array[43849] = 16'h12d7;
mem_array[43848] = 16'h3d69;
mem_array[43851] = 16'h07d2;
mem_array[43850] = 16'h3d2b;
mem_array[43853] = 16'h1259;
mem_array[43852] = 16'hbd79;
mem_array[43855] = 16'h23ff;
mem_array[43854] = 16'h3cc4;
mem_array[43857] = 16'hde58;
mem_array[43856] = 16'hbd8c;
mem_array[43859] = 16'hd288;
mem_array[43858] = 16'hbcbf;
mem_array[43861] = 16'ha917;
mem_array[43860] = 16'h3d90;
mem_array[43863] = 16'h399a;
mem_array[43862] = 16'h3d3b;
mem_array[43865] = 16'h2b8f;
mem_array[43864] = 16'h3db1;
mem_array[43867] = 16'h1867;
mem_array[43866] = 16'h3d1a;
mem_array[43869] = 16'h6e0f;
mem_array[43868] = 16'hbc0f;
mem_array[43871] = 16'h2863;
mem_array[43870] = 16'h3d2e;
mem_array[43873] = 16'haaa1;
mem_array[43872] = 16'h3c42;
mem_array[43875] = 16'h42dd;
mem_array[43874] = 16'h3c89;
mem_array[43877] = 16'hc3f3;
mem_array[43876] = 16'h3c48;
mem_array[43879] = 16'h4b2b;
mem_array[43878] = 16'hbd99;
mem_array[43881] = 16'hb957;
mem_array[43880] = 16'h3cb1;
mem_array[43883] = 16'h0e6f;
mem_array[43882] = 16'hbd3e;
mem_array[43885] = 16'h239a;
mem_array[43884] = 16'h3ca6;
mem_array[43887] = 16'hea6f;
mem_array[43886] = 16'h3b78;
mem_array[43889] = 16'h6a1e;
mem_array[43888] = 16'hbd6e;
mem_array[43891] = 16'h6574;
mem_array[43890] = 16'hbd07;
mem_array[43893] = 16'h9329;
mem_array[43892] = 16'hbd43;
mem_array[43895] = 16'hd282;
mem_array[43894] = 16'hbc46;
mem_array[43897] = 16'h05da;
mem_array[43896] = 16'h3cbf;
mem_array[43899] = 16'h0ce3;
mem_array[43898] = 16'h3c23;
mem_array[43901] = 16'hf4c0;
mem_array[43900] = 16'h3da3;
mem_array[43903] = 16'h784c;
mem_array[43902] = 16'h3d63;
mem_array[43905] = 16'hf438;
mem_array[43904] = 16'h3dcb;
mem_array[43907] = 16'h1ca4;
mem_array[43906] = 16'hbc75;
mem_array[43909] = 16'h3333;
mem_array[43908] = 16'hbbed;
mem_array[43911] = 16'hb5f8;
mem_array[43910] = 16'h3db8;
mem_array[43913] = 16'h1dfe;
mem_array[43912] = 16'hbd0c;
mem_array[43915] = 16'hc708;
mem_array[43914] = 16'hbd3c;
mem_array[43917] = 16'h343e;
mem_array[43916] = 16'h3ca5;
mem_array[43919] = 16'hc4ba;
mem_array[43918] = 16'hbd9d;
mem_array[43921] = 16'hc7c3;
mem_array[43920] = 16'hbd13;
mem_array[43923] = 16'h8c57;
mem_array[43922] = 16'h3f2a;
mem_array[43925] = 16'h9159;
mem_array[43924] = 16'hbf44;
mem_array[43927] = 16'hbe61;
mem_array[43926] = 16'h3cde;
mem_array[43929] = 16'h970b;
mem_array[43928] = 16'h3ee8;
mem_array[43931] = 16'hd3e7;
mem_array[43930] = 16'hbeab;
mem_array[43933] = 16'hfef5;
mem_array[43932] = 16'hbf1c;
mem_array[43935] = 16'h02a6;
mem_array[43934] = 16'hbf24;
mem_array[43937] = 16'h719f;
mem_array[43936] = 16'h38ac;
mem_array[43939] = 16'h80d0;
mem_array[43938] = 16'hbddc;
mem_array[43941] = 16'hfdc1;
mem_array[43940] = 16'h3d08;
mem_array[43943] = 16'h20ca;
mem_array[43942] = 16'hbd79;
mem_array[43945] = 16'hd73b;
mem_array[43944] = 16'hbda1;
mem_array[43947] = 16'he423;
mem_array[43946] = 16'hbd8f;
mem_array[43949] = 16'hd5ef;
mem_array[43948] = 16'h3e5e;
mem_array[43951] = 16'h2ee5;
mem_array[43950] = 16'h3f08;
mem_array[43953] = 16'h3d88;
mem_array[43952] = 16'hbe40;
mem_array[43955] = 16'h6455;
mem_array[43954] = 16'hbeb9;
mem_array[43957] = 16'h3f2e;
mem_array[43956] = 16'h3e0b;
mem_array[43959] = 16'h8fdc;
mem_array[43958] = 16'h3e23;
mem_array[43961] = 16'h1a7e;
mem_array[43960] = 16'h3dc9;
mem_array[43963] = 16'h0442;
mem_array[43962] = 16'hbf19;
mem_array[43965] = 16'hdc9d;
mem_array[43964] = 16'h3d0f;
mem_array[43967] = 16'h3447;
mem_array[43966] = 16'h3f2c;
mem_array[43969] = 16'h2706;
mem_array[43968] = 16'hbed5;
mem_array[43971] = 16'h04e2;
mem_array[43970] = 16'hbef4;
mem_array[43973] = 16'h04dd;
mem_array[43972] = 16'hbe87;
mem_array[43975] = 16'h03f7;
mem_array[43974] = 16'h3d2f;
mem_array[43977] = 16'hfc97;
mem_array[43976] = 16'hbdba;
mem_array[43979] = 16'hb39e;
mem_array[43978] = 16'h3e97;
mem_array[43981] = 16'h153a;
mem_array[43980] = 16'hbe32;
mem_array[43983] = 16'heeaf;
mem_array[43982] = 16'hbea1;
mem_array[43985] = 16'h6e03;
mem_array[43984] = 16'hbf0f;
mem_array[43987] = 16'h51fc;
mem_array[43986] = 16'hbea2;
mem_array[43989] = 16'h8c07;
mem_array[43988] = 16'h3edc;
mem_array[43991] = 16'hca56;
mem_array[43990] = 16'hbf31;
mem_array[43993] = 16'he74e;
mem_array[43992] = 16'hbf04;
mem_array[43995] = 16'h8db2;
mem_array[43994] = 16'h3e93;
mem_array[43997] = 16'h56e0;
mem_array[43996] = 16'h3c95;
mem_array[43999] = 16'hd987;
mem_array[43998] = 16'h3c19;
mem_array[44001] = 16'h41fb;
mem_array[44000] = 16'h3cd4;
mem_array[44003] = 16'h8f2d;
mem_array[44002] = 16'hbdb6;
mem_array[44005] = 16'h894d;
mem_array[44004] = 16'hbec0;
mem_array[44007] = 16'ha5b3;
mem_array[44006] = 16'hbdf4;
mem_array[44009] = 16'hb915;
mem_array[44008] = 16'h3eed;
mem_array[44011] = 16'h576d;
mem_array[44010] = 16'h3db1;
mem_array[44013] = 16'h2001;
mem_array[44012] = 16'hbebc;
mem_array[44015] = 16'hef1d;
mem_array[44014] = 16'hbf07;
mem_array[44017] = 16'h0f00;
mem_array[44016] = 16'hbf4e;
mem_array[44019] = 16'h4e51;
mem_array[44018] = 16'h3df9;
mem_array[44021] = 16'h057d;
mem_array[44020] = 16'hbefe;
mem_array[44023] = 16'h3d98;
mem_array[44022] = 16'hbf00;
mem_array[44025] = 16'h0c0e;
mem_array[44024] = 16'hbd35;
mem_array[44027] = 16'h1c59;
mem_array[44026] = 16'h3f6c;
mem_array[44029] = 16'h2026;
mem_array[44028] = 16'h3d67;
mem_array[44031] = 16'h3c1f;
mem_array[44030] = 16'hbfab;
mem_array[44033] = 16'h342b;
mem_array[44032] = 16'hbf03;
mem_array[44035] = 16'h98e3;
mem_array[44034] = 16'hbe67;
mem_array[44037] = 16'h4f8e;
mem_array[44036] = 16'hbe2e;
mem_array[44039] = 16'h3eff;
mem_array[44038] = 16'h3e58;
mem_array[44041] = 16'hbcc2;
mem_array[44040] = 16'hbecc;
mem_array[44043] = 16'h8bd7;
mem_array[44042] = 16'hbe60;
mem_array[44045] = 16'h9621;
mem_array[44044] = 16'hbec9;
mem_array[44047] = 16'hf35a;
mem_array[44046] = 16'hbea6;
mem_array[44049] = 16'hff63;
mem_array[44048] = 16'h3ecb;
mem_array[44051] = 16'hd063;
mem_array[44050] = 16'hbe24;
mem_array[44053] = 16'h9c4d;
mem_array[44052] = 16'hbeac;
mem_array[44055] = 16'h292d;
mem_array[44054] = 16'h3f3b;
mem_array[44057] = 16'hdb07;
mem_array[44056] = 16'hbecd;
mem_array[44059] = 16'h2172;
mem_array[44058] = 16'h3e43;
mem_array[44061] = 16'h6c06;
mem_array[44060] = 16'hbd00;
mem_array[44063] = 16'h0ff9;
mem_array[44062] = 16'hbd02;
mem_array[44065] = 16'h1b01;
mem_array[44064] = 16'hbf1c;
mem_array[44067] = 16'h7799;
mem_array[44066] = 16'hbc83;
mem_array[44069] = 16'hc24f;
mem_array[44068] = 16'h3ea8;
mem_array[44071] = 16'h6a0b;
mem_array[44070] = 16'hbe64;
mem_array[44073] = 16'h2d4f;
mem_array[44072] = 16'hbe02;
mem_array[44075] = 16'hcf45;
mem_array[44074] = 16'h3d48;
mem_array[44077] = 16'h448b;
mem_array[44076] = 16'hbedd;
mem_array[44079] = 16'h24e8;
mem_array[44078] = 16'h3e57;
mem_array[44081] = 16'h1865;
mem_array[44080] = 16'hbf0c;
mem_array[44083] = 16'hc2d5;
mem_array[44082] = 16'hbe88;
mem_array[44085] = 16'h1f5b;
mem_array[44084] = 16'h3d67;
mem_array[44087] = 16'h50f3;
mem_array[44086] = 16'h3e52;
mem_array[44089] = 16'hfd36;
mem_array[44088] = 16'hbd8d;
mem_array[44091] = 16'he0c2;
mem_array[44090] = 16'hbf3c;
mem_array[44093] = 16'h5288;
mem_array[44092] = 16'hbed0;
mem_array[44095] = 16'h6895;
mem_array[44094] = 16'hbeb5;
mem_array[44097] = 16'hfe2d;
mem_array[44096] = 16'hbd85;
mem_array[44099] = 16'h3c65;
mem_array[44098] = 16'h3e05;
mem_array[44101] = 16'ha588;
mem_array[44100] = 16'hbf57;
mem_array[44103] = 16'h5ca9;
mem_array[44102] = 16'h3e23;
mem_array[44105] = 16'h0539;
mem_array[44104] = 16'hbd32;
mem_array[44107] = 16'hde85;
mem_array[44106] = 16'hbe52;
mem_array[44109] = 16'ha8e5;
mem_array[44108] = 16'h3f3e;
mem_array[44111] = 16'h2354;
mem_array[44110] = 16'h3f3b;
mem_array[44113] = 16'h667d;
mem_array[44112] = 16'hbf81;
mem_array[44115] = 16'h0adf;
mem_array[44114] = 16'h3f6d;
mem_array[44117] = 16'ha43e;
mem_array[44116] = 16'h3ea3;
mem_array[44119] = 16'h24c0;
mem_array[44118] = 16'h3e58;
mem_array[44121] = 16'hec75;
mem_array[44120] = 16'h3c6b;
mem_array[44123] = 16'h20a4;
mem_array[44122] = 16'h3c32;
mem_array[44125] = 16'h94be;
mem_array[44124] = 16'hbff2;
mem_array[44127] = 16'h3277;
mem_array[44126] = 16'h3d94;
mem_array[44129] = 16'he042;
mem_array[44128] = 16'h3eb0;
mem_array[44131] = 16'hf87c;
mem_array[44130] = 16'hbdec;
mem_array[44133] = 16'h29a0;
mem_array[44132] = 16'hbec7;
mem_array[44135] = 16'h7b36;
mem_array[44134] = 16'h3e5c;
mem_array[44137] = 16'h5697;
mem_array[44136] = 16'h3eb1;
mem_array[44139] = 16'ha3a2;
mem_array[44138] = 16'hbc4b;
mem_array[44141] = 16'h418b;
mem_array[44140] = 16'hbfac;
mem_array[44143] = 16'h0b71;
mem_array[44142] = 16'h3ec7;
mem_array[44145] = 16'hc1f2;
mem_array[44144] = 16'h3c26;
mem_array[44147] = 16'h8a28;
mem_array[44146] = 16'hbe9a;
mem_array[44149] = 16'h1eb4;
mem_array[44148] = 16'h3c7c;
mem_array[44151] = 16'h5f18;
mem_array[44150] = 16'h3f3e;
mem_array[44153] = 16'h4bf3;
mem_array[44152] = 16'h3eae;
mem_array[44155] = 16'he486;
mem_array[44154] = 16'hbe66;
mem_array[44157] = 16'hec1f;
mem_array[44156] = 16'h3d38;
mem_array[44159] = 16'h5c9c;
mem_array[44158] = 16'hbec5;
mem_array[44161] = 16'h14f2;
mem_array[44160] = 16'hbf80;
mem_array[44163] = 16'h5666;
mem_array[44162] = 16'h3ea2;
mem_array[44165] = 16'hd121;
mem_array[44164] = 16'h3e0c;
mem_array[44167] = 16'hbdc4;
mem_array[44166] = 16'hbefa;
mem_array[44169] = 16'h9ccf;
mem_array[44168] = 16'hbd96;
mem_array[44171] = 16'h2810;
mem_array[44170] = 16'hbebe;
mem_array[44173] = 16'hcb7b;
mem_array[44172] = 16'h3c91;
mem_array[44175] = 16'h91d9;
mem_array[44174] = 16'h3ed5;
mem_array[44177] = 16'h5add;
mem_array[44176] = 16'h3e50;
mem_array[44179] = 16'hfc8a;
mem_array[44178] = 16'h3e9b;
mem_array[44181] = 16'h6d24;
mem_array[44180] = 16'hbd08;
mem_array[44183] = 16'h73a6;
mem_array[44182] = 16'hbda5;
mem_array[44185] = 16'hbedb;
mem_array[44184] = 16'hbfa5;
mem_array[44187] = 16'h7634;
mem_array[44186] = 16'hbe3b;
mem_array[44189] = 16'h9272;
mem_array[44188] = 16'h3f47;
mem_array[44191] = 16'h0289;
mem_array[44190] = 16'h3e28;
mem_array[44193] = 16'h0505;
mem_array[44192] = 16'hbf83;
mem_array[44195] = 16'h31fb;
mem_array[44194] = 16'h3f6f;
mem_array[44197] = 16'hb6f4;
mem_array[44196] = 16'h3ed2;
mem_array[44199] = 16'ha8a4;
mem_array[44198] = 16'hbef9;
mem_array[44201] = 16'h8376;
mem_array[44200] = 16'hbf3e;
mem_array[44203] = 16'hf3b9;
mem_array[44202] = 16'h3ea9;
mem_array[44205] = 16'h8ba0;
mem_array[44204] = 16'h3c4c;
mem_array[44207] = 16'h3a7e;
mem_array[44206] = 16'h3e36;
mem_array[44209] = 16'h785e;
mem_array[44208] = 16'h3ee4;
mem_array[44211] = 16'h5e84;
mem_array[44210] = 16'h3f33;
mem_array[44213] = 16'h1944;
mem_array[44212] = 16'h3e83;
mem_array[44215] = 16'h7c7c;
mem_array[44214] = 16'hbf5a;
mem_array[44217] = 16'hb1ae;
mem_array[44216] = 16'hbe87;
mem_array[44219] = 16'hce4e;
mem_array[44218] = 16'hbf6e;
mem_array[44221] = 16'haadf;
mem_array[44220] = 16'hbed4;
mem_array[44223] = 16'hab49;
mem_array[44222] = 16'h3ecd;
mem_array[44225] = 16'hb368;
mem_array[44224] = 16'h3ea8;
mem_array[44227] = 16'hccea;
mem_array[44226] = 16'hbfa7;
mem_array[44229] = 16'hf1fc;
mem_array[44228] = 16'hbeaa;
mem_array[44231] = 16'hdf5c;
mem_array[44230] = 16'hbf01;
mem_array[44233] = 16'h799f;
mem_array[44232] = 16'h3e24;
mem_array[44235] = 16'hac75;
mem_array[44234] = 16'hbe95;
mem_array[44237] = 16'he9ff;
mem_array[44236] = 16'hbf6b;
mem_array[44239] = 16'h2b33;
mem_array[44238] = 16'hbdfd;
mem_array[44241] = 16'h8cb1;
mem_array[44240] = 16'h3d38;
mem_array[44243] = 16'habe2;
mem_array[44242] = 16'h3ca2;
mem_array[44245] = 16'hbcc9;
mem_array[44244] = 16'hbf11;
mem_array[44247] = 16'ha7f0;
mem_array[44246] = 16'hbf0a;
mem_array[44249] = 16'h653e;
mem_array[44248] = 16'h3ee3;
mem_array[44251] = 16'hc5a5;
mem_array[44250] = 16'h3e84;
mem_array[44253] = 16'he395;
mem_array[44252] = 16'hbf3b;
mem_array[44255] = 16'h858b;
mem_array[44254] = 16'h3d04;
mem_array[44257] = 16'hfdd2;
mem_array[44256] = 16'h3fa8;
mem_array[44259] = 16'ha8bb;
mem_array[44258] = 16'hbf8d;
mem_array[44261] = 16'hcbc6;
mem_array[44260] = 16'hbf78;
mem_array[44263] = 16'hc8cb;
mem_array[44262] = 16'h3f01;
mem_array[44265] = 16'h0c27;
mem_array[44264] = 16'h3dc5;
mem_array[44267] = 16'h6b53;
mem_array[44266] = 16'h3f09;
mem_array[44269] = 16'h6871;
mem_array[44268] = 16'hbe7b;
mem_array[44271] = 16'he95f;
mem_array[44270] = 16'hbe18;
mem_array[44273] = 16'h91a8;
mem_array[44272] = 16'h3e14;
mem_array[44275] = 16'hf2a0;
mem_array[44274] = 16'hbe91;
mem_array[44277] = 16'h87e3;
mem_array[44276] = 16'hbeed;
mem_array[44279] = 16'had34;
mem_array[44278] = 16'hbfdc;
mem_array[44281] = 16'h7152;
mem_array[44280] = 16'hbe86;
mem_array[44283] = 16'h3f1b;
mem_array[44282] = 16'h3c10;
mem_array[44285] = 16'h033d;
mem_array[44284] = 16'h3f15;
mem_array[44287] = 16'hd73c;
mem_array[44286] = 16'hbfa1;
mem_array[44289] = 16'hf0a6;
mem_array[44288] = 16'h3f26;
mem_array[44291] = 16'hd2a4;
mem_array[44290] = 16'h3f01;
mem_array[44293] = 16'h460a;
mem_array[44292] = 16'hbd70;
mem_array[44295] = 16'hebf4;
mem_array[44294] = 16'hbe4a;
mem_array[44297] = 16'hb764;
mem_array[44296] = 16'hbf4b;
mem_array[44299] = 16'hf674;
mem_array[44298] = 16'h3d72;
mem_array[44301] = 16'hf1ca;
mem_array[44300] = 16'h3c20;
mem_array[44303] = 16'ha904;
mem_array[44302] = 16'h3d80;
mem_array[44305] = 16'hfa51;
mem_array[44304] = 16'hbf06;
mem_array[44307] = 16'ha648;
mem_array[44306] = 16'hbeba;
mem_array[44309] = 16'h8d00;
mem_array[44308] = 16'h3eb6;
mem_array[44311] = 16'hd987;
mem_array[44310] = 16'h3e11;
mem_array[44313] = 16'h9345;
mem_array[44312] = 16'hbe3e;
mem_array[44315] = 16'hc5f7;
mem_array[44314] = 16'hbe94;
mem_array[44317] = 16'h0665;
mem_array[44316] = 16'h3ef8;
mem_array[44319] = 16'heddd;
mem_array[44318] = 16'hbe91;
mem_array[44321] = 16'hf38f;
mem_array[44320] = 16'hbf3a;
mem_array[44323] = 16'h5e39;
mem_array[44322] = 16'h3f1e;
mem_array[44325] = 16'h9c6f;
mem_array[44324] = 16'h3e9e;
mem_array[44327] = 16'h046b;
mem_array[44326] = 16'h3ece;
mem_array[44329] = 16'hd935;
mem_array[44328] = 16'h3eac;
mem_array[44331] = 16'hf830;
mem_array[44330] = 16'hbf55;
mem_array[44333] = 16'hc36f;
mem_array[44332] = 16'h3e13;
mem_array[44335] = 16'hda8a;
mem_array[44334] = 16'hbeb6;
mem_array[44337] = 16'h0067;
mem_array[44336] = 16'hbd8f;
mem_array[44339] = 16'h8e42;
mem_array[44338] = 16'hbfc5;
mem_array[44341] = 16'h4ba9;
mem_array[44340] = 16'hbea3;
mem_array[44343] = 16'he257;
mem_array[44342] = 16'h3db6;
mem_array[44345] = 16'h924f;
mem_array[44344] = 16'h3c34;
mem_array[44347] = 16'h0317;
mem_array[44346] = 16'hbefa;
mem_array[44349] = 16'h909f;
mem_array[44348] = 16'h3f84;
mem_array[44351] = 16'h17d0;
mem_array[44350] = 16'h3edf;
mem_array[44353] = 16'h198c;
mem_array[44352] = 16'hbe49;
mem_array[44355] = 16'h7bfa;
mem_array[44354] = 16'h3f10;
mem_array[44357] = 16'h6548;
mem_array[44356] = 16'h3e32;
mem_array[44359] = 16'h0bbf;
mem_array[44358] = 16'hbf01;
mem_array[44361] = 16'hf6ca;
mem_array[44360] = 16'h3bf3;
mem_array[44363] = 16'h727f;
mem_array[44362] = 16'hbda2;
mem_array[44365] = 16'h2bd2;
mem_array[44364] = 16'hbf0d;
mem_array[44367] = 16'h6976;
mem_array[44366] = 16'hbf0a;
mem_array[44369] = 16'hfc7c;
mem_array[44368] = 16'hbf3a;
mem_array[44371] = 16'h1f09;
mem_array[44370] = 16'hbdb7;
mem_array[44373] = 16'h9e2b;
mem_array[44372] = 16'hbf3a;
mem_array[44375] = 16'h8e51;
mem_array[44374] = 16'hbf81;
mem_array[44377] = 16'hb189;
mem_array[44376] = 16'h3b9c;
mem_array[44379] = 16'hea07;
mem_array[44378] = 16'hbe11;
mem_array[44381] = 16'h4c59;
mem_array[44380] = 16'hbf0a;
mem_array[44383] = 16'h3db7;
mem_array[44382] = 16'h3f0b;
mem_array[44385] = 16'h367e;
mem_array[44384] = 16'h3e10;
mem_array[44387] = 16'haf55;
mem_array[44386] = 16'h3f1b;
mem_array[44389] = 16'h3f92;
mem_array[44388] = 16'h3ee0;
mem_array[44391] = 16'hf6d6;
mem_array[44390] = 16'hbf4a;
mem_array[44393] = 16'hf654;
mem_array[44392] = 16'h3f25;
mem_array[44395] = 16'heb46;
mem_array[44394] = 16'hbe98;
mem_array[44397] = 16'hef3a;
mem_array[44396] = 16'hbe97;
mem_array[44399] = 16'h9dee;
mem_array[44398] = 16'hbf68;
mem_array[44401] = 16'h6294;
mem_array[44400] = 16'hbf57;
mem_array[44403] = 16'hd033;
mem_array[44402] = 16'hbe09;
mem_array[44405] = 16'hd3e1;
mem_array[44404] = 16'hbe8d;
mem_array[44407] = 16'h8254;
mem_array[44406] = 16'hbf0d;
mem_array[44409] = 16'hb7c1;
mem_array[44408] = 16'h3e50;
mem_array[44411] = 16'had97;
mem_array[44410] = 16'hbf24;
mem_array[44413] = 16'hdf2d;
mem_array[44412] = 16'h3e30;
mem_array[44415] = 16'h595d;
mem_array[44414] = 16'h3f40;
mem_array[44417] = 16'h8f5f;
mem_array[44416] = 16'h3e2b;
mem_array[44419] = 16'hac49;
mem_array[44418] = 16'hbfa5;
mem_array[44421] = 16'he018;
mem_array[44420] = 16'hbd83;
mem_array[44423] = 16'h510b;
mem_array[44422] = 16'hbd96;
mem_array[44425] = 16'hbe68;
mem_array[44424] = 16'hbefe;
mem_array[44427] = 16'h097e;
mem_array[44426] = 16'hbe75;
mem_array[44429] = 16'h78af;
mem_array[44428] = 16'hbea1;
mem_array[44431] = 16'h04f5;
mem_array[44430] = 16'hbe49;
mem_array[44433] = 16'hf752;
mem_array[44432] = 16'hbf32;
mem_array[44435] = 16'hee7c;
mem_array[44434] = 16'hbee2;
mem_array[44437] = 16'h9569;
mem_array[44436] = 16'h3ea4;
mem_array[44439] = 16'he9b5;
mem_array[44438] = 16'h3d76;
mem_array[44441] = 16'hcc68;
mem_array[44440] = 16'hbf66;
mem_array[44443] = 16'hd50f;
mem_array[44442] = 16'h3f24;
mem_array[44445] = 16'hfa81;
mem_array[44444] = 16'h3e18;
mem_array[44447] = 16'hee07;
mem_array[44446] = 16'h3ef7;
mem_array[44449] = 16'hc9c4;
mem_array[44448] = 16'hbe07;
mem_array[44451] = 16'h464e;
mem_array[44450] = 16'hbf19;
mem_array[44453] = 16'h7cf2;
mem_array[44452] = 16'h3ec6;
mem_array[44455] = 16'ha9a4;
mem_array[44454] = 16'h3d40;
mem_array[44457] = 16'hd10a;
mem_array[44456] = 16'hbdbf;
mem_array[44459] = 16'hda1e;
mem_array[44458] = 16'hc01b;
mem_array[44461] = 16'hf977;
mem_array[44460] = 16'h3f38;
mem_array[44463] = 16'h2bd1;
mem_array[44462] = 16'h3eb8;
mem_array[44465] = 16'hbb6a;
mem_array[44464] = 16'h3f5c;
mem_array[44467] = 16'h4021;
mem_array[44466] = 16'hbfb7;
mem_array[44469] = 16'h0eb8;
mem_array[44468] = 16'h3ef9;
mem_array[44471] = 16'h63a7;
mem_array[44470] = 16'h3ee8;
mem_array[44473] = 16'he2e5;
mem_array[44472] = 16'h3f08;
mem_array[44475] = 16'h6856;
mem_array[44474] = 16'h3f14;
mem_array[44477] = 16'h0a60;
mem_array[44476] = 16'hbdaa;
mem_array[44479] = 16'h3495;
mem_array[44478] = 16'hbf34;
mem_array[44481] = 16'hd376;
mem_array[44480] = 16'hbd1b;
mem_array[44483] = 16'h40eb;
mem_array[44482] = 16'h39bb;
mem_array[44485] = 16'ha76a;
mem_array[44484] = 16'hbfa9;
mem_array[44487] = 16'hc7b1;
mem_array[44486] = 16'hbdeb;
mem_array[44489] = 16'h471a;
mem_array[44488] = 16'hbeac;
mem_array[44491] = 16'hc06c;
mem_array[44490] = 16'hbe66;
mem_array[44493] = 16'hab65;
mem_array[44492] = 16'hbde9;
mem_array[44495] = 16'hb704;
mem_array[44494] = 16'hbf04;
mem_array[44497] = 16'h5e53;
mem_array[44496] = 16'h3ecb;
mem_array[44499] = 16'hd91e;
mem_array[44498] = 16'hbe26;
mem_array[44501] = 16'ha993;
mem_array[44500] = 16'hbf6d;
mem_array[44503] = 16'h3976;
mem_array[44502] = 16'h3f14;
mem_array[44505] = 16'h59a8;
mem_array[44504] = 16'h3dcf;
mem_array[44507] = 16'hc286;
mem_array[44506] = 16'h3f14;
mem_array[44509] = 16'he8b6;
mem_array[44508] = 16'hbd83;
mem_array[44511] = 16'h693d;
mem_array[44510] = 16'h3eb0;
mem_array[44513] = 16'h14af;
mem_array[44512] = 16'h3f1f;
mem_array[44515] = 16'h18f9;
mem_array[44514] = 16'h3f28;
mem_array[44517] = 16'h0b68;
mem_array[44516] = 16'h3f12;
mem_array[44519] = 16'h9c4f;
mem_array[44518] = 16'hbf16;
mem_array[44521] = 16'h4360;
mem_array[44520] = 16'hbc8b;
mem_array[44523] = 16'h4f51;
mem_array[44522] = 16'h3e84;
mem_array[44525] = 16'h1f5a;
mem_array[44524] = 16'h3f1d;
mem_array[44527] = 16'h5a77;
mem_array[44526] = 16'hbf81;
mem_array[44529] = 16'hb060;
mem_array[44528] = 16'h3eb2;
mem_array[44531] = 16'hf8cd;
mem_array[44530] = 16'hbec6;
mem_array[44533] = 16'h3156;
mem_array[44532] = 16'hbf71;
mem_array[44535] = 16'hf336;
mem_array[44534] = 16'h3daa;
mem_array[44537] = 16'h3a32;
mem_array[44536] = 16'hbefd;
mem_array[44539] = 16'ha424;
mem_array[44538] = 16'hbf9d;
mem_array[44541] = 16'hf47a;
mem_array[44540] = 16'hbd7f;
mem_array[44543] = 16'h38e6;
mem_array[44542] = 16'h3d48;
mem_array[44545] = 16'hb9e8;
mem_array[44544] = 16'hbf98;
mem_array[44547] = 16'h61b4;
mem_array[44546] = 16'hbecb;
mem_array[44549] = 16'hffd1;
mem_array[44548] = 16'h3e9c;
mem_array[44551] = 16'h63e5;
mem_array[44550] = 16'h3ed5;
mem_array[44553] = 16'hb412;
mem_array[44552] = 16'hbecb;
mem_array[44555] = 16'h4525;
mem_array[44554] = 16'hbf28;
mem_array[44557] = 16'hc2c6;
mem_array[44556] = 16'h3f10;
mem_array[44559] = 16'h3c7f;
mem_array[44558] = 16'hbf59;
mem_array[44561] = 16'hd689;
mem_array[44560] = 16'hbf7b;
mem_array[44563] = 16'hc032;
mem_array[44562] = 16'h3e8f;
mem_array[44565] = 16'h3ce2;
mem_array[44564] = 16'hbda2;
mem_array[44567] = 16'h0c81;
mem_array[44566] = 16'h3ef7;
mem_array[44569] = 16'h91b2;
mem_array[44568] = 16'h3edf;
mem_array[44571] = 16'h4eb1;
mem_array[44570] = 16'h3c78;
mem_array[44573] = 16'hb34c;
mem_array[44572] = 16'h3e90;
mem_array[44575] = 16'h5df2;
mem_array[44574] = 16'hbebb;
mem_array[44577] = 16'hb7c2;
mem_array[44576] = 16'h3e38;
mem_array[44579] = 16'hd5e1;
mem_array[44578] = 16'hbf25;
mem_array[44581] = 16'h2540;
mem_array[44580] = 16'hbeea;
mem_array[44583] = 16'h483a;
mem_array[44582] = 16'h3e9d;
mem_array[44585] = 16'h89c5;
mem_array[44584] = 16'h3e93;
mem_array[44587] = 16'h7d02;
mem_array[44586] = 16'hbf83;
mem_array[44589] = 16'hb6a9;
mem_array[44588] = 16'h3ec7;
mem_array[44591] = 16'hdbed;
mem_array[44590] = 16'hbdb7;
mem_array[44593] = 16'hf459;
mem_array[44592] = 16'hbf9a;
mem_array[44595] = 16'hcc27;
mem_array[44594] = 16'hbd57;
mem_array[44597] = 16'h6e47;
mem_array[44596] = 16'hbf9f;
mem_array[44599] = 16'h8108;
mem_array[44598] = 16'hbf33;
mem_array[44601] = 16'hf7f5;
mem_array[44600] = 16'h3b54;
mem_array[44603] = 16'h19bd;
mem_array[44602] = 16'hbd87;
mem_array[44605] = 16'h4a77;
mem_array[44604] = 16'hbe71;
mem_array[44607] = 16'hec94;
mem_array[44606] = 16'hbef0;
mem_array[44609] = 16'hc542;
mem_array[44608] = 16'hbe41;
mem_array[44611] = 16'h3f60;
mem_array[44610] = 16'h3c3f;
mem_array[44613] = 16'h5398;
mem_array[44612] = 16'hbda7;
mem_array[44615] = 16'h0c5d;
mem_array[44614] = 16'hbfab;
mem_array[44617] = 16'h27c2;
mem_array[44616] = 16'h3d7f;
mem_array[44619] = 16'h085b;
mem_array[44618] = 16'hbed8;
mem_array[44621] = 16'h5258;
mem_array[44620] = 16'hbf8d;
mem_array[44623] = 16'hc66c;
mem_array[44622] = 16'h3ee4;
mem_array[44625] = 16'h9e4f;
mem_array[44624] = 16'h3e7a;
mem_array[44627] = 16'h479a;
mem_array[44626] = 16'h3f7d;
mem_array[44629] = 16'he8f2;
mem_array[44628] = 16'hbd5c;
mem_array[44631] = 16'h94b4;
mem_array[44630] = 16'hbe92;
mem_array[44633] = 16'h8732;
mem_array[44632] = 16'h3f05;
mem_array[44635] = 16'ha4af;
mem_array[44634] = 16'hbeee;
mem_array[44637] = 16'h9c05;
mem_array[44636] = 16'h3eb9;
mem_array[44639] = 16'h16ce;
mem_array[44638] = 16'h3c01;
mem_array[44641] = 16'h238f;
mem_array[44640] = 16'h3f14;
mem_array[44643] = 16'hd198;
mem_array[44642] = 16'h3e72;
mem_array[44645] = 16'hae29;
mem_array[44644] = 16'h3dfb;
mem_array[44647] = 16'hed43;
mem_array[44646] = 16'hbf5b;
mem_array[44649] = 16'h4ccf;
mem_array[44648] = 16'h3e66;
mem_array[44651] = 16'h1573;
mem_array[44650] = 16'hbee5;
mem_array[44653] = 16'h94ff;
mem_array[44652] = 16'hbf36;
mem_array[44655] = 16'h1fc0;
mem_array[44654] = 16'h3e9a;
mem_array[44657] = 16'he454;
mem_array[44656] = 16'h3e81;
mem_array[44659] = 16'hc8fc;
mem_array[44658] = 16'h3e31;
mem_array[44661] = 16'h075e;
mem_array[44660] = 16'hbd1a;
mem_array[44663] = 16'h7a65;
mem_array[44662] = 16'h3c68;
mem_array[44665] = 16'hc122;
mem_array[44664] = 16'hbf4d;
mem_array[44667] = 16'h4da5;
mem_array[44666] = 16'hbe41;
mem_array[44669] = 16'h1b90;
mem_array[44668] = 16'hbf7c;
mem_array[44671] = 16'hcd24;
mem_array[44670] = 16'hbe20;
mem_array[44673] = 16'h4b91;
mem_array[44672] = 16'hbea6;
mem_array[44675] = 16'hc6d5;
mem_array[44674] = 16'hbf41;
mem_array[44677] = 16'h4203;
mem_array[44676] = 16'h3e95;
mem_array[44679] = 16'hda55;
mem_array[44678] = 16'hbe88;
mem_array[44681] = 16'h2fc3;
mem_array[44680] = 16'hbf8f;
mem_array[44683] = 16'hd710;
mem_array[44682] = 16'hbcb3;
mem_array[44685] = 16'h11ed;
mem_array[44684] = 16'h3e26;
mem_array[44687] = 16'h22b9;
mem_array[44686] = 16'h3e89;
mem_array[44689] = 16'hc67b;
mem_array[44688] = 16'h3e16;
mem_array[44691] = 16'ha388;
mem_array[44690] = 16'h3e8e;
mem_array[44693] = 16'h16a4;
mem_array[44692] = 16'hbdcf;
mem_array[44695] = 16'h8acc;
mem_array[44694] = 16'h3f02;
mem_array[44697] = 16'h73f3;
mem_array[44696] = 16'h3f09;
mem_array[44699] = 16'hf0c2;
mem_array[44698] = 16'hbf53;
mem_array[44701] = 16'hbae8;
mem_array[44700] = 16'h3edc;
mem_array[44703] = 16'haf64;
mem_array[44702] = 16'h3bf3;
mem_array[44705] = 16'h4096;
mem_array[44704] = 16'hbf00;
mem_array[44707] = 16'hf12e;
mem_array[44706] = 16'hbfca;
mem_array[44709] = 16'hb237;
mem_array[44708] = 16'hbec8;
mem_array[44711] = 16'ha082;
mem_array[44710] = 16'hbf6f;
mem_array[44713] = 16'h0957;
mem_array[44712] = 16'h3f07;
mem_array[44715] = 16'h1d5f;
mem_array[44714] = 16'h3dad;
mem_array[44717] = 16'hb03a;
mem_array[44716] = 16'hbed5;
mem_array[44719] = 16'h1fc2;
mem_array[44718] = 16'hbee5;
mem_array[44721] = 16'h3a61;
mem_array[44720] = 16'hbda3;
mem_array[44723] = 16'h5f51;
mem_array[44722] = 16'h3ceb;
mem_array[44725] = 16'hec78;
mem_array[44724] = 16'hbf0e;
mem_array[44727] = 16'hca00;
mem_array[44726] = 16'hbd85;
mem_array[44729] = 16'hdbb9;
mem_array[44728] = 16'hbf81;
mem_array[44731] = 16'h4f1f;
mem_array[44730] = 16'h3e72;
mem_array[44733] = 16'h3186;
mem_array[44732] = 16'hbedd;
mem_array[44735] = 16'h81b8;
mem_array[44734] = 16'hbf67;
mem_array[44737] = 16'hcc47;
mem_array[44736] = 16'h3e40;
mem_array[44739] = 16'hc610;
mem_array[44738] = 16'hbe7a;
mem_array[44741] = 16'h0a90;
mem_array[44740] = 16'hbfa1;
mem_array[44743] = 16'hce01;
mem_array[44742] = 16'hbe03;
mem_array[44745] = 16'hbab4;
mem_array[44744] = 16'h3dad;
mem_array[44747] = 16'h36ac;
mem_array[44746] = 16'h3efe;
mem_array[44749] = 16'h5fed;
mem_array[44748] = 16'hbe7e;
mem_array[44751] = 16'h91cc;
mem_array[44750] = 16'h3de9;
mem_array[44753] = 16'h2230;
mem_array[44752] = 16'hbe61;
mem_array[44755] = 16'h869e;
mem_array[44754] = 16'h3ebe;
mem_array[44757] = 16'hbe0f;
mem_array[44756] = 16'h3f07;
mem_array[44759] = 16'hc555;
mem_array[44758] = 16'hbf4d;
mem_array[44761] = 16'h1af1;
mem_array[44760] = 16'h3ebc;
mem_array[44763] = 16'hee19;
mem_array[44762] = 16'hbe6f;
mem_array[44765] = 16'h1f97;
mem_array[44764] = 16'h3ddf;
mem_array[44767] = 16'hbab1;
mem_array[44766] = 16'hbfb4;
mem_array[44769] = 16'h1da2;
mem_array[44768] = 16'h3d18;
mem_array[44771] = 16'h72d1;
mem_array[44770] = 16'hbf1f;
mem_array[44773] = 16'hb411;
mem_array[44772] = 16'h3f2e;
mem_array[44775] = 16'h8679;
mem_array[44774] = 16'h3e19;
mem_array[44777] = 16'hf13c;
mem_array[44776] = 16'hbe8c;
mem_array[44779] = 16'hb4a4;
mem_array[44778] = 16'hbe13;
mem_array[44781] = 16'h1da7;
mem_array[44780] = 16'hbd80;
mem_array[44783] = 16'hbfa3;
mem_array[44782] = 16'hbd6e;
mem_array[44785] = 16'hd5f1;
mem_array[44784] = 16'hbf31;
mem_array[44787] = 16'h626c;
mem_array[44786] = 16'hbe1c;
mem_array[44789] = 16'h0a10;
mem_array[44788] = 16'hbf81;
mem_array[44791] = 16'h1b2e;
mem_array[44790] = 16'hbe3a;
mem_array[44793] = 16'hf982;
mem_array[44792] = 16'hbed8;
mem_array[44795] = 16'h7638;
mem_array[44794] = 16'hbfa8;
mem_array[44797] = 16'hffee;
mem_array[44796] = 16'h3e1f;
mem_array[44799] = 16'hfc6d;
mem_array[44798] = 16'hbf8b;
mem_array[44801] = 16'h8b52;
mem_array[44800] = 16'hbf34;
mem_array[44803] = 16'hdf47;
mem_array[44802] = 16'hbd2b;
mem_array[44805] = 16'h2e4a;
mem_array[44804] = 16'h3d27;
mem_array[44807] = 16'h2cae;
mem_array[44806] = 16'h3f0d;
mem_array[44809] = 16'h9e2c;
mem_array[44808] = 16'h3e4b;
mem_array[44811] = 16'h8b14;
mem_array[44810] = 16'h3f82;
mem_array[44813] = 16'hf64a;
mem_array[44812] = 16'h3e75;
mem_array[44815] = 16'h0f3d;
mem_array[44814] = 16'h3e60;
mem_array[44817] = 16'h033b;
mem_array[44816] = 16'h3e50;
mem_array[44819] = 16'h29e8;
mem_array[44818] = 16'hbfc1;
mem_array[44821] = 16'hda78;
mem_array[44820] = 16'h3ea2;
mem_array[44823] = 16'hce1d;
mem_array[44822] = 16'h3fbd;
mem_array[44825] = 16'hc7e2;
mem_array[44824] = 16'h3f30;
mem_array[44827] = 16'hc46c;
mem_array[44826] = 16'h3ea4;
mem_array[44829] = 16'h67d9;
mem_array[44828] = 16'hbf9a;
mem_array[44831] = 16'hd457;
mem_array[44830] = 16'h3ecc;
mem_array[44833] = 16'hbbfc;
mem_array[44832] = 16'h3f0e;
mem_array[44835] = 16'h821c;
mem_array[44834] = 16'h3d64;
mem_array[44837] = 16'he867;
mem_array[44836] = 16'hbe82;
mem_array[44839] = 16'hdcbc;
mem_array[44838] = 16'hbe55;
mem_array[44841] = 16'h6129;
mem_array[44840] = 16'hbd3d;
mem_array[44843] = 16'h3a66;
mem_array[44842] = 16'h3bd7;
mem_array[44845] = 16'h4d50;
mem_array[44844] = 16'hbe6e;
mem_array[44847] = 16'hfea4;
mem_array[44846] = 16'hbe4f;
mem_array[44849] = 16'h2a4d;
mem_array[44848] = 16'hbd3f;
mem_array[44851] = 16'hec6a;
mem_array[44850] = 16'hbf21;
mem_array[44853] = 16'h5e56;
mem_array[44852] = 16'h3d36;
mem_array[44855] = 16'h1e65;
mem_array[44854] = 16'hbf2c;
mem_array[44857] = 16'h8636;
mem_array[44856] = 16'hbd94;
mem_array[44859] = 16'h78bb;
mem_array[44858] = 16'hbf74;
mem_array[44861] = 16'h8027;
mem_array[44860] = 16'hbf8a;
mem_array[44863] = 16'h8ae7;
mem_array[44862] = 16'hbe86;
mem_array[44865] = 16'h1960;
mem_array[44864] = 16'h3de7;
mem_array[44867] = 16'hb452;
mem_array[44866] = 16'h3e2f;
mem_array[44869] = 16'h8f4e;
mem_array[44868] = 16'h3cf7;
mem_array[44871] = 16'hda2e;
mem_array[44870] = 16'h3f6a;
mem_array[44873] = 16'ha16d;
mem_array[44872] = 16'h3e9f;
mem_array[44875] = 16'he5b1;
mem_array[44874] = 16'h3e9d;
mem_array[44877] = 16'ha690;
mem_array[44876] = 16'hbeb5;
mem_array[44879] = 16'h41f3;
mem_array[44878] = 16'hc008;
mem_array[44881] = 16'h9e80;
mem_array[44880] = 16'hbc5b;
mem_array[44883] = 16'he872;
mem_array[44882] = 16'hbf07;
mem_array[44885] = 16'h0620;
mem_array[44884] = 16'hbde6;
mem_array[44887] = 16'h6c9e;
mem_array[44886] = 16'hbf71;
mem_array[44889] = 16'h32b2;
mem_array[44888] = 16'h3ea4;
mem_array[44891] = 16'hd794;
mem_array[44890] = 16'h3e0e;
mem_array[44893] = 16'hbfc6;
mem_array[44892] = 16'h3f82;
mem_array[44895] = 16'hd9bd;
mem_array[44894] = 16'hbe54;
mem_array[44897] = 16'h902c;
mem_array[44896] = 16'hbe60;
mem_array[44899] = 16'h97af;
mem_array[44898] = 16'hbefc;
mem_array[44901] = 16'h8464;
mem_array[44900] = 16'hbd70;
mem_array[44903] = 16'ha1ca;
mem_array[44902] = 16'hbcdb;
mem_array[44905] = 16'h366e;
mem_array[44904] = 16'hbe3b;
mem_array[44907] = 16'h9f8c;
mem_array[44906] = 16'hbe20;
mem_array[44909] = 16'h1504;
mem_array[44908] = 16'hbf03;
mem_array[44911] = 16'hf3ba;
mem_array[44910] = 16'h3eb8;
mem_array[44913] = 16'h3a08;
mem_array[44912] = 16'hbdfa;
mem_array[44915] = 16'h3368;
mem_array[44914] = 16'hbf60;
mem_array[44917] = 16'h679f;
mem_array[44916] = 16'h3e2c;
mem_array[44919] = 16'hc224;
mem_array[44918] = 16'hbe03;
mem_array[44921] = 16'hcdd6;
mem_array[44920] = 16'hbf9e;
mem_array[44923] = 16'h652a;
mem_array[44922] = 16'hbe32;
mem_array[44925] = 16'h5cf4;
mem_array[44924] = 16'h3b04;
mem_array[44927] = 16'h03fe;
mem_array[44926] = 16'hbe95;
mem_array[44929] = 16'h9976;
mem_array[44928] = 16'hbf02;
mem_array[44931] = 16'h139f;
mem_array[44930] = 16'hbe61;
mem_array[44933] = 16'h1dd3;
mem_array[44932] = 16'h3ec3;
mem_array[44935] = 16'hc16e;
mem_array[44934] = 16'hbeb9;
mem_array[44937] = 16'hdf78;
mem_array[44936] = 16'hbf16;
mem_array[44939] = 16'h6dea;
mem_array[44938] = 16'hc007;
mem_array[44941] = 16'h51b3;
mem_array[44940] = 16'hbce0;
mem_array[44943] = 16'h9c50;
mem_array[44942] = 16'hbe81;
mem_array[44945] = 16'h3658;
mem_array[44944] = 16'hbf89;
mem_array[44947] = 16'hc4b0;
mem_array[44946] = 16'hbf24;
mem_array[44949] = 16'h1b09;
mem_array[44948] = 16'h3f5c;
mem_array[44951] = 16'hdb8a;
mem_array[44950] = 16'h3d11;
mem_array[44953] = 16'h32a0;
mem_array[44952] = 16'h3f25;
mem_array[44955] = 16'h4f0b;
mem_array[44954] = 16'h3f5d;
mem_array[44957] = 16'ha616;
mem_array[44956] = 16'hbf2e;
mem_array[44959] = 16'h323a;
mem_array[44958] = 16'hbd24;
mem_array[44961] = 16'h3dcc;
mem_array[44960] = 16'hbd51;
mem_array[44963] = 16'h65b9;
mem_array[44962] = 16'hbdc3;
mem_array[44965] = 16'h602a;
mem_array[44964] = 16'hbf2e;
mem_array[44967] = 16'ha623;
mem_array[44966] = 16'hbdaf;
mem_array[44969] = 16'hddf5;
mem_array[44968] = 16'hbe48;
mem_array[44971] = 16'h7d24;
mem_array[44970] = 16'h3e88;
mem_array[44973] = 16'h287b;
mem_array[44972] = 16'hbdbf;
mem_array[44975] = 16'h5531;
mem_array[44974] = 16'hbfb9;
mem_array[44977] = 16'h6ff1;
mem_array[44976] = 16'h3f19;
mem_array[44979] = 16'h4b92;
mem_array[44978] = 16'hbf2e;
mem_array[44981] = 16'h1ac7;
mem_array[44980] = 16'hbfd8;
mem_array[44983] = 16'hbcc0;
mem_array[44982] = 16'h3e9f;
mem_array[44985] = 16'haef4;
mem_array[44984] = 16'h3beb;
mem_array[44987] = 16'h1b4d;
mem_array[44986] = 16'hbf20;
mem_array[44989] = 16'h8a53;
mem_array[44988] = 16'hbf31;
mem_array[44991] = 16'hac5f;
mem_array[44990] = 16'h3dc3;
mem_array[44993] = 16'h7607;
mem_array[44992] = 16'h3e45;
mem_array[44995] = 16'h1a61;
mem_array[44994] = 16'h3f43;
mem_array[44997] = 16'h2b33;
mem_array[44996] = 16'hbda2;
mem_array[44999] = 16'hf7bb;
mem_array[44998] = 16'hbfb1;
mem_array[45001] = 16'h05f4;
mem_array[45000] = 16'h3cab;
mem_array[45003] = 16'h9a17;
mem_array[45002] = 16'h3e82;
mem_array[45005] = 16'hf976;
mem_array[45004] = 16'hbec2;
mem_array[45007] = 16'hdb11;
mem_array[45006] = 16'h3d93;
mem_array[45009] = 16'h97e8;
mem_array[45008] = 16'h3ef0;
mem_array[45011] = 16'h3395;
mem_array[45010] = 16'hbd72;
mem_array[45013] = 16'h27f8;
mem_array[45012] = 16'h3f50;
mem_array[45015] = 16'h7138;
mem_array[45014] = 16'h3f59;
mem_array[45017] = 16'h977d;
mem_array[45016] = 16'hbe5a;
mem_array[45019] = 16'ha10a;
mem_array[45018] = 16'h3cf1;
mem_array[45021] = 16'hc1e8;
mem_array[45020] = 16'hbcb1;
mem_array[45023] = 16'h2da6;
mem_array[45022] = 16'hbc13;
mem_array[45025] = 16'h4b67;
mem_array[45024] = 16'h3e7b;
mem_array[45027] = 16'h9dcf;
mem_array[45026] = 16'hbea5;
mem_array[45029] = 16'h9adb;
mem_array[45028] = 16'hbe47;
mem_array[45031] = 16'h639b;
mem_array[45030] = 16'hbf00;
mem_array[45033] = 16'hfa04;
mem_array[45032] = 16'hbd90;
mem_array[45035] = 16'h9aec;
mem_array[45034] = 16'hbf87;
mem_array[45037] = 16'h4d76;
mem_array[45036] = 16'hbd28;
mem_array[45039] = 16'h3abc;
mem_array[45038] = 16'hbf90;
mem_array[45041] = 16'hc0b5;
mem_array[45040] = 16'hbfd0;
mem_array[45043] = 16'hfe80;
mem_array[45042] = 16'h3f23;
mem_array[45045] = 16'he701;
mem_array[45044] = 16'hbcd4;
mem_array[45047] = 16'hb056;
mem_array[45046] = 16'hbcb2;
mem_array[45049] = 16'ha88f;
mem_array[45048] = 16'hbdf1;
mem_array[45051] = 16'hbbca;
mem_array[45050] = 16'h3ef9;
mem_array[45053] = 16'h8600;
mem_array[45052] = 16'h3f12;
mem_array[45055] = 16'h582b;
mem_array[45054] = 16'h3ea3;
mem_array[45057] = 16'hc398;
mem_array[45056] = 16'hbca2;
mem_array[45059] = 16'hf93a;
mem_array[45058] = 16'hbf6f;
mem_array[45061] = 16'h8d6a;
mem_array[45060] = 16'hbdaa;
mem_array[45063] = 16'h2f2a;
mem_array[45062] = 16'h3f89;
mem_array[45065] = 16'hd73a;
mem_array[45064] = 16'h3c9a;
mem_array[45067] = 16'h9065;
mem_array[45066] = 16'h3e18;
mem_array[45069] = 16'h016b;
mem_array[45068] = 16'hbf4e;
mem_array[45071] = 16'hd8a7;
mem_array[45070] = 16'hbded;
mem_array[45073] = 16'ha8ff;
mem_array[45072] = 16'h3b92;
mem_array[45075] = 16'h03eb;
mem_array[45074] = 16'h3f25;
mem_array[45077] = 16'h3946;
mem_array[45076] = 16'h3acd;
mem_array[45079] = 16'h350d;
mem_array[45078] = 16'hbda3;
mem_array[45081] = 16'hada0;
mem_array[45080] = 16'h3d81;
mem_array[45083] = 16'h47e8;
mem_array[45082] = 16'h3d38;
mem_array[45085] = 16'h2f35;
mem_array[45084] = 16'h3e7f;
mem_array[45087] = 16'he010;
mem_array[45086] = 16'h3c7e;
mem_array[45089] = 16'hb552;
mem_array[45088] = 16'h3de2;
mem_array[45091] = 16'hc15e;
mem_array[45090] = 16'h3b9f;
mem_array[45093] = 16'hfd5b;
mem_array[45092] = 16'hbbd8;
mem_array[45095] = 16'hd2b2;
mem_array[45094] = 16'hbf3b;
mem_array[45097] = 16'h9eaf;
mem_array[45096] = 16'h3efc;
mem_array[45099] = 16'hce8c;
mem_array[45098] = 16'hbe23;
mem_array[45101] = 16'h3c53;
mem_array[45100] = 16'hbf82;
mem_array[45103] = 16'ha393;
mem_array[45102] = 16'hbdc5;
mem_array[45105] = 16'h178c;
mem_array[45104] = 16'hbd40;
mem_array[45107] = 16'h1e07;
mem_array[45106] = 16'hbe56;
mem_array[45109] = 16'h6c26;
mem_array[45108] = 16'hbda3;
mem_array[45111] = 16'h1907;
mem_array[45110] = 16'h3ebe;
mem_array[45113] = 16'h7df5;
mem_array[45112] = 16'h3f0f;
mem_array[45115] = 16'h746f;
mem_array[45114] = 16'h3f0f;
mem_array[45117] = 16'h3c9c;
mem_array[45116] = 16'hbd58;
mem_array[45119] = 16'h8862;
mem_array[45118] = 16'hbf24;
mem_array[45121] = 16'h7cd8;
mem_array[45120] = 16'h3c77;
mem_array[45123] = 16'hec17;
mem_array[45122] = 16'hbe78;
mem_array[45125] = 16'hde7e;
mem_array[45124] = 16'hbc74;
mem_array[45127] = 16'he9bd;
mem_array[45126] = 16'hbbaa;
mem_array[45129] = 16'h8cae;
mem_array[45128] = 16'h3e86;
mem_array[45131] = 16'h682c;
mem_array[45130] = 16'h3b81;
mem_array[45133] = 16'ha5e6;
mem_array[45132] = 16'hbcc8;
mem_array[45135] = 16'h1e80;
mem_array[45134] = 16'hbdb0;
mem_array[45137] = 16'hc6e6;
mem_array[45136] = 16'h3de9;
mem_array[45139] = 16'hd180;
mem_array[45138] = 16'hbd04;
mem_array[45141] = 16'h127f;
mem_array[45140] = 16'hbd38;
mem_array[45143] = 16'h0601;
mem_array[45142] = 16'hbdbe;
mem_array[45145] = 16'hd967;
mem_array[45144] = 16'h3ea8;
mem_array[45147] = 16'h4dbb;
mem_array[45146] = 16'h3d5f;
mem_array[45149] = 16'h1f0a;
mem_array[45148] = 16'hbd26;
mem_array[45151] = 16'h36b8;
mem_array[45150] = 16'h3f2a;
mem_array[45153] = 16'h37d8;
mem_array[45152] = 16'h3c09;
mem_array[45155] = 16'hfb64;
mem_array[45154] = 16'hbd42;
mem_array[45157] = 16'h3233;
mem_array[45156] = 16'h3f23;
mem_array[45159] = 16'hf0b8;
mem_array[45158] = 16'h3e92;
mem_array[45161] = 16'h2f66;
mem_array[45160] = 16'h3e24;
mem_array[45163] = 16'h3ded;
mem_array[45162] = 16'hbeef;
mem_array[45165] = 16'h551c;
mem_array[45164] = 16'hbce1;
mem_array[45167] = 16'hd5ee;
mem_array[45166] = 16'hbf1e;
mem_array[45169] = 16'h71f7;
mem_array[45168] = 16'h3dd1;
mem_array[45171] = 16'ha37d;
mem_array[45170] = 16'hbec4;
mem_array[45173] = 16'hdb51;
mem_array[45172] = 16'hbca9;
mem_array[45175] = 16'h6ae9;
mem_array[45174] = 16'h3d1b;
mem_array[45177] = 16'h9554;
mem_array[45176] = 16'h3b82;
mem_array[45179] = 16'hf3c8;
mem_array[45178] = 16'hbe0b;
mem_array[45181] = 16'h21d0;
mem_array[45180] = 16'hbdb8;
mem_array[45183] = 16'h3bb3;
mem_array[45182] = 16'hbda7;
mem_array[45185] = 16'h4e8d;
mem_array[45184] = 16'h3d8a;
mem_array[45187] = 16'hf4d3;
mem_array[45186] = 16'hbd8a;
mem_array[45189] = 16'h7204;
mem_array[45188] = 16'h3bf0;
mem_array[45191] = 16'hdadd;
mem_array[45190] = 16'hbe2d;
mem_array[45193] = 16'h3813;
mem_array[45192] = 16'hbdaf;
mem_array[45195] = 16'h70bf;
mem_array[45194] = 16'hbd45;
mem_array[45197] = 16'h6206;
mem_array[45196] = 16'hbcbe;
mem_array[45199] = 16'he289;
mem_array[45198] = 16'h3c84;
mem_array[45201] = 16'hfacd;
mem_array[45200] = 16'h3b07;
mem_array[45203] = 16'h7034;
mem_array[45202] = 16'hbcad;
mem_array[45205] = 16'h183e;
mem_array[45204] = 16'h3d01;
mem_array[45207] = 16'h6214;
mem_array[45206] = 16'hbd23;
mem_array[45209] = 16'he00e;
mem_array[45208] = 16'hbd03;
mem_array[45211] = 16'hb3d2;
mem_array[45210] = 16'h3ca6;
mem_array[45213] = 16'h632e;
mem_array[45212] = 16'h3bdb;
mem_array[45215] = 16'h4562;
mem_array[45214] = 16'hbdb4;
mem_array[45217] = 16'hebfa;
mem_array[45216] = 16'h3d90;
mem_array[45219] = 16'hd23e;
mem_array[45218] = 16'hbd7c;
mem_array[45221] = 16'h5499;
mem_array[45220] = 16'h3b6b;
mem_array[45223] = 16'he193;
mem_array[45222] = 16'h3d87;
mem_array[45225] = 16'hd896;
mem_array[45224] = 16'h3da1;
mem_array[45227] = 16'h658c;
mem_array[45226] = 16'hbc84;
mem_array[45229] = 16'h4914;
mem_array[45228] = 16'hbd6c;
mem_array[45231] = 16'h2e7f;
mem_array[45230] = 16'h3c4a;
mem_array[45233] = 16'h6a68;
mem_array[45232] = 16'hbb97;
mem_array[45235] = 16'hfd0a;
mem_array[45234] = 16'h3dd4;
mem_array[45237] = 16'h8a38;
mem_array[45236] = 16'h3c1e;
mem_array[45239] = 16'h7563;
mem_array[45238] = 16'hbc30;
mem_array[45241] = 16'h708f;
mem_array[45240] = 16'h3c3f;
mem_array[45243] = 16'h9a2a;
mem_array[45242] = 16'h3ce9;
mem_array[45245] = 16'h799b;
mem_array[45244] = 16'h3c37;
mem_array[45247] = 16'h0ac8;
mem_array[45246] = 16'hbdeb;
mem_array[45249] = 16'h1940;
mem_array[45248] = 16'h3d0f;
mem_array[45251] = 16'ha36c;
mem_array[45250] = 16'hbd09;
mem_array[45253] = 16'h8126;
mem_array[45252] = 16'h3d57;
mem_array[45255] = 16'h0074;
mem_array[45254] = 16'h3cc0;
mem_array[45257] = 16'hb8dd;
mem_array[45256] = 16'hbb2a;
mem_array[45259] = 16'hb2a5;
mem_array[45258] = 16'h3cb9;
mem_array[45261] = 16'h45f9;
mem_array[45260] = 16'hba42;
mem_array[45263] = 16'hdb8d;
mem_array[45262] = 16'h3d76;
mem_array[45265] = 16'ha077;
mem_array[45264] = 16'hbda8;
mem_array[45267] = 16'he40c;
mem_array[45266] = 16'hbca3;
mem_array[45269] = 16'h9553;
mem_array[45268] = 16'h3d04;
mem_array[45271] = 16'h9e16;
mem_array[45270] = 16'h3ce1;
mem_array[45273] = 16'h6b84;
mem_array[45272] = 16'hbd1c;
mem_array[45275] = 16'h6239;
mem_array[45274] = 16'hbd1c;
mem_array[45277] = 16'h9af5;
mem_array[45276] = 16'h3cb5;
mem_array[45279] = 16'h9cfc;
mem_array[45278] = 16'h3d0a;
mem_array[45281] = 16'hced6;
mem_array[45280] = 16'hbc2f;
mem_array[45283] = 16'h70c0;
mem_array[45282] = 16'hbd8d;
mem_array[45285] = 16'h6013;
mem_array[45284] = 16'hbdd8;
mem_array[45287] = 16'hb9a8;
mem_array[45286] = 16'h3d77;
mem_array[45289] = 16'h2569;
mem_array[45288] = 16'hbd36;
mem_array[45291] = 16'haccc;
mem_array[45290] = 16'hbd1e;
mem_array[45293] = 16'h6d66;
mem_array[45292] = 16'hbd8e;
mem_array[45295] = 16'hea58;
mem_array[45294] = 16'hbcca;
mem_array[45297] = 16'h8ead;
mem_array[45296] = 16'hbd67;
mem_array[45299] = 16'h3ba3;
mem_array[45298] = 16'hbb2f;
mem_array[45301] = 16'h4cea;
mem_array[45300] = 16'h3b24;
mem_array[45303] = 16'h277c;
mem_array[45302] = 16'h3bb0;
mem_array[45305] = 16'h3ad4;
mem_array[45304] = 16'h3d3c;
mem_array[45307] = 16'h341d;
mem_array[45306] = 16'h3c09;
mem_array[45309] = 16'h08f8;
mem_array[45308] = 16'hbcd3;
mem_array[45311] = 16'h090d;
mem_array[45310] = 16'hbd32;
mem_array[45313] = 16'ha3a4;
mem_array[45312] = 16'hb978;
mem_array[45315] = 16'h8edd;
mem_array[45314] = 16'hbc2f;
mem_array[45317] = 16'h78d3;
mem_array[45316] = 16'h3d31;
mem_array[45319] = 16'h669a;
mem_array[45318] = 16'h3ce9;
mem_array[45321] = 16'hfe55;
mem_array[45320] = 16'h3d1f;
mem_array[45323] = 16'ha4ba;
mem_array[45322] = 16'hbc87;
mem_array[45325] = 16'hd986;
mem_array[45324] = 16'h3d93;
mem_array[45327] = 16'hadca;
mem_array[45326] = 16'h3d38;
mem_array[45329] = 16'h9bdb;
mem_array[45328] = 16'h3ca0;
mem_array[45331] = 16'h924f;
mem_array[45330] = 16'hbb90;
mem_array[45333] = 16'h74e8;
mem_array[45332] = 16'h3caf;
mem_array[45335] = 16'head2;
mem_array[45334] = 16'hbd38;
mem_array[45337] = 16'hda74;
mem_array[45336] = 16'h3d95;
mem_array[45339] = 16'hd143;
mem_array[45338] = 16'hbcbb;
mem_array[45341] = 16'h3940;
mem_array[45340] = 16'h3c7c;
mem_array[45343] = 16'h728d;
mem_array[45342] = 16'hbc5d;
mem_array[45345] = 16'h0775;
mem_array[45344] = 16'hbd3d;
mem_array[45347] = 16'hd96f;
mem_array[45346] = 16'h3d01;
mem_array[45349] = 16'h230f;
mem_array[45348] = 16'hbd66;
mem_array[45351] = 16'h0581;
mem_array[45350] = 16'h3c8e;
mem_array[45353] = 16'h1ea3;
mem_array[45352] = 16'hbcc1;
mem_array[45355] = 16'h6d63;
mem_array[45354] = 16'h3d10;
mem_array[45357] = 16'h05dc;
mem_array[45356] = 16'hbd81;
mem_array[45359] = 16'hc006;
mem_array[45358] = 16'hbd65;
mem_array[45361] = 16'h53d6;
mem_array[45360] = 16'hbd97;
mem_array[45363] = 16'h6f6e;
mem_array[45362] = 16'h3d84;
mem_array[45365] = 16'hfde7;
mem_array[45364] = 16'hbd46;
mem_array[45367] = 16'hda3f;
mem_array[45366] = 16'h3dbf;
mem_array[45369] = 16'h7619;
mem_array[45368] = 16'h3d28;
mem_array[45371] = 16'h636b;
mem_array[45370] = 16'h3dcc;
mem_array[45373] = 16'h4c69;
mem_array[45372] = 16'hbcd6;
mem_array[45375] = 16'h5c7b;
mem_array[45374] = 16'h3b93;
mem_array[45377] = 16'h2d29;
mem_array[45376] = 16'hbda4;
mem_array[45379] = 16'ha213;
mem_array[45378] = 16'hbce2;
mem_array[45381] = 16'h9023;
mem_array[45380] = 16'hbd1f;
mem_array[45383] = 16'h92de;
mem_array[45382] = 16'h3d20;
mem_array[45385] = 16'h3104;
mem_array[45384] = 16'hbdc3;
mem_array[45387] = 16'hefdb;
mem_array[45386] = 16'hbd40;
mem_array[45389] = 16'he8c5;
mem_array[45388] = 16'hbd57;
mem_array[45391] = 16'h369f;
mem_array[45390] = 16'hbca8;
mem_array[45393] = 16'h1e68;
mem_array[45392] = 16'h3d26;
mem_array[45395] = 16'hf911;
mem_array[45394] = 16'h3d49;
mem_array[45397] = 16'h5843;
mem_array[45396] = 16'h3b5e;
mem_array[45399] = 16'hbe15;
mem_array[45398] = 16'h3cff;
mem_array[45401] = 16'h57d6;
mem_array[45400] = 16'hbd37;
mem_array[45403] = 16'ha540;
mem_array[45402] = 16'h3d36;
mem_array[45405] = 16'h831d;
mem_array[45404] = 16'hbcf8;
mem_array[45407] = 16'hd650;
mem_array[45406] = 16'h3db4;
mem_array[45409] = 16'h9acc;
mem_array[45408] = 16'hbd84;
mem_array[45411] = 16'h6895;
mem_array[45410] = 16'hbda9;
mem_array[45413] = 16'hb14a;
mem_array[45412] = 16'hbc12;
mem_array[45415] = 16'hda24;
mem_array[45414] = 16'h3d5b;
mem_array[45417] = 16'h78c4;
mem_array[45416] = 16'hbbec;
mem_array[45419] = 16'h660b;
mem_array[45418] = 16'hbbd8;
mem_array[45421] = 16'h7297;
mem_array[45420] = 16'h3d49;
mem_array[45423] = 16'h3637;
mem_array[45422] = 16'hbd39;
mem_array[45425] = 16'h4f0f;
mem_array[45424] = 16'hbc2b;
mem_array[45427] = 16'hdd4b;
mem_array[45426] = 16'h3daa;
mem_array[45429] = 16'h5da3;
mem_array[45428] = 16'hbcc9;
mem_array[45431] = 16'hfeb4;
mem_array[45430] = 16'hbd7d;
mem_array[45433] = 16'h83fd;
mem_array[45432] = 16'h3c40;
mem_array[45435] = 16'h6d59;
mem_array[45434] = 16'hbc52;
mem_array[45437] = 16'h4fa4;
mem_array[45436] = 16'h3d81;
mem_array[45439] = 16'h2275;
mem_array[45438] = 16'hbda5;
mem_array[45441] = 16'h5aaa;
mem_array[45440] = 16'h3d05;
mem_array[45443] = 16'h5664;
mem_array[45442] = 16'h3d78;
mem_array[45445] = 16'h7156;
mem_array[45444] = 16'hbd16;
mem_array[45447] = 16'h2431;
mem_array[45446] = 16'h3d46;
mem_array[45449] = 16'haa48;
mem_array[45448] = 16'h3ce2;
mem_array[45451] = 16'h66fa;
mem_array[45450] = 16'hbc03;
mem_array[45453] = 16'h53f6;
mem_array[45452] = 16'h3d4d;
mem_array[45455] = 16'h465a;
mem_array[45454] = 16'hbde1;
mem_array[45457] = 16'h2eb1;
mem_array[45456] = 16'h3c7f;
mem_array[45459] = 16'h27ac;
mem_array[45458] = 16'h3cc6;
mem_array[45461] = 16'hc6d0;
mem_array[45460] = 16'h3dc2;
mem_array[45463] = 16'h85cb;
mem_array[45462] = 16'h3dda;
mem_array[45465] = 16'hb456;
mem_array[45464] = 16'h3ddc;
mem_array[45467] = 16'h7660;
mem_array[45466] = 16'h3d3a;
mem_array[45469] = 16'h7be4;
mem_array[45468] = 16'h3d87;
mem_array[45471] = 16'hfc10;
mem_array[45470] = 16'h3be4;
mem_array[45473] = 16'h064f;
mem_array[45472] = 16'hbd1e;
mem_array[45475] = 16'h2938;
mem_array[45474] = 16'h3db7;
mem_array[45477] = 16'hfad5;
mem_array[45476] = 16'hbd78;
mem_array[45479] = 16'h9c7f;
mem_array[45478] = 16'h3da5;
mem_array[45481] = 16'h016d;
mem_array[45480] = 16'hbca2;
mem_array[45483] = 16'h5aed;
mem_array[45482] = 16'hbd86;
mem_array[45485] = 16'h193b;
mem_array[45484] = 16'hbc59;
mem_array[45487] = 16'hb8c5;
mem_array[45486] = 16'hbd39;
mem_array[45489] = 16'h87fd;
mem_array[45488] = 16'hbccf;
mem_array[45491] = 16'h90d0;
mem_array[45490] = 16'hbde0;
mem_array[45493] = 16'hca6c;
mem_array[45492] = 16'h3db1;
mem_array[45495] = 16'ha364;
mem_array[45494] = 16'h3ca7;
mem_array[45497] = 16'hb043;
mem_array[45496] = 16'h3d57;
mem_array[45499] = 16'h4be9;
mem_array[45498] = 16'h3cd5;
mem_array[45501] = 16'he566;
mem_array[45500] = 16'h3dce;
mem_array[45503] = 16'hd3c6;
mem_array[45502] = 16'hbd48;
mem_array[45505] = 16'hf223;
mem_array[45504] = 16'h3d2a;
mem_array[45507] = 16'hf5a2;
mem_array[45506] = 16'hbdab;
mem_array[45509] = 16'h2992;
mem_array[45508] = 16'h3ccc;
mem_array[45511] = 16'hcb22;
mem_array[45510] = 16'hbc9f;
mem_array[45513] = 16'hac84;
mem_array[45512] = 16'hbd84;
mem_array[45515] = 16'h5a2d;
mem_array[45514] = 16'hbd54;
mem_array[45517] = 16'hb556;
mem_array[45516] = 16'h3da2;
mem_array[45519] = 16'hbbf3;
mem_array[45518] = 16'hbbc7;
mem_array[45521] = 16'h375c;
mem_array[45520] = 16'h3c62;
mem_array[45523] = 16'h3f05;
mem_array[45522] = 16'h3c9f;
mem_array[45525] = 16'h5eaa;
mem_array[45524] = 16'hbd07;
mem_array[45527] = 16'h0200;
mem_array[45526] = 16'hbc30;
mem_array[45529] = 16'h9500;
mem_array[45528] = 16'h3d19;
mem_array[45531] = 16'hbd7d;
mem_array[45530] = 16'hbda2;
mem_array[45533] = 16'h0176;
mem_array[45532] = 16'hbca6;
mem_array[45535] = 16'hf6a3;
mem_array[45534] = 16'hbd22;
mem_array[45537] = 16'h5d9d;
mem_array[45536] = 16'hbb19;
mem_array[45539] = 16'hc94f;
mem_array[45538] = 16'h3c6d;
mem_array[45541] = 16'hcef9;
mem_array[45540] = 16'hbcfb;
mem_array[45543] = 16'h1c56;
mem_array[45542] = 16'hbddc;
mem_array[45545] = 16'he9cd;
mem_array[45544] = 16'h3dea;
mem_array[45547] = 16'hcf06;
mem_array[45546] = 16'hbd50;
mem_array[45549] = 16'h3d53;
mem_array[45548] = 16'hbdbc;
mem_array[45551] = 16'h1369;
mem_array[45550] = 16'hbcee;
mem_array[45553] = 16'hf874;
mem_array[45552] = 16'h3cdd;
mem_array[45555] = 16'h46eb;
mem_array[45554] = 16'h3d19;
mem_array[45557] = 16'hf272;
mem_array[45556] = 16'h3d8b;
mem_array[45559] = 16'h558b;
mem_array[45558] = 16'hbcad;
mem_array[45561] = 16'hc2f5;
mem_array[45560] = 16'hbd22;
mem_array[45563] = 16'h8dc0;
mem_array[45562] = 16'h3c67;
mem_array[45565] = 16'he11e;
mem_array[45564] = 16'h3c0b;
mem_array[45567] = 16'h5ec6;
mem_array[45566] = 16'h3d97;
mem_array[45569] = 16'hac8f;
mem_array[45568] = 16'h3c8d;
mem_array[45571] = 16'h31b3;
mem_array[45570] = 16'hbd92;
mem_array[45573] = 16'h3a94;
mem_array[45572] = 16'hbce6;
mem_array[45575] = 16'hdb34;
mem_array[45574] = 16'h3d2f;
mem_array[45577] = 16'h5246;
mem_array[45576] = 16'h3dae;
mem_array[45579] = 16'h261d;
mem_array[45578] = 16'hbd07;
mem_array[45581] = 16'hb7b3;
mem_array[45580] = 16'hbbc4;
mem_array[45583] = 16'h42b0;
mem_array[45582] = 16'h3d27;
mem_array[45585] = 16'hd551;
mem_array[45584] = 16'h3d3c;
mem_array[45587] = 16'hac90;
mem_array[45586] = 16'h3c73;
mem_array[45589] = 16'ha33e;
mem_array[45588] = 16'h3cd6;
mem_array[45591] = 16'h6d20;
mem_array[45590] = 16'hbdcf;
mem_array[45593] = 16'h8bb6;
mem_array[45592] = 16'hbc99;
mem_array[45595] = 16'h2e84;
mem_array[45594] = 16'hbce0;
mem_array[45597] = 16'h61e8;
mem_array[45596] = 16'hbd2f;
mem_array[45599] = 16'h03b4;
mem_array[45598] = 16'hb924;
mem_array[45601] = 16'hbb40;
mem_array[45600] = 16'hbd90;
mem_array[45603] = 16'h71cd;
mem_array[45602] = 16'h3d53;
mem_array[45605] = 16'he0b8;
mem_array[45604] = 16'h3e06;
mem_array[45607] = 16'h9202;
mem_array[45606] = 16'h3d59;
mem_array[45609] = 16'h1948;
mem_array[45608] = 16'h3edd;
mem_array[45611] = 16'h0f83;
mem_array[45610] = 16'hbe14;
mem_array[45613] = 16'h9853;
mem_array[45612] = 16'h3d3f;
mem_array[45615] = 16'hce2b;
mem_array[45614] = 16'h3d62;
mem_array[45617] = 16'he983;
mem_array[45616] = 16'h3dd4;
mem_array[45619] = 16'h6a42;
mem_array[45618] = 16'h3c80;
mem_array[45621] = 16'hd4f9;
mem_array[45620] = 16'hbd2f;
mem_array[45623] = 16'he813;
mem_array[45622] = 16'h3d09;
mem_array[45625] = 16'hd9cb;
mem_array[45624] = 16'h3d9e;
mem_array[45627] = 16'hfda4;
mem_array[45626] = 16'h3d83;
mem_array[45629] = 16'hfdb0;
mem_array[45628] = 16'h3e44;
mem_array[45631] = 16'h7fd8;
mem_array[45630] = 16'hbe98;
mem_array[45633] = 16'h316c;
mem_array[45632] = 16'h3bc2;
mem_array[45635] = 16'hb307;
mem_array[45634] = 16'hbcd6;
mem_array[45637] = 16'ha2ef;
mem_array[45636] = 16'h3e15;
mem_array[45639] = 16'ha1f3;
mem_array[45638] = 16'h3d13;
mem_array[45641] = 16'h6cf0;
mem_array[45640] = 16'hbc82;
mem_array[45643] = 16'hdec4;
mem_array[45642] = 16'hbe52;
mem_array[45645] = 16'h07e3;
mem_array[45644] = 16'h3d51;
mem_array[45647] = 16'hff6e;
mem_array[45646] = 16'hbf3d;
mem_array[45649] = 16'h857c;
mem_array[45648] = 16'hbb94;
mem_array[45651] = 16'hb11b;
mem_array[45650] = 16'h3f4c;
mem_array[45653] = 16'h9508;
mem_array[45652] = 16'hbe2e;
mem_array[45655] = 16'hf273;
mem_array[45654] = 16'h3e9f;
mem_array[45657] = 16'hb08a;
mem_array[45656] = 16'h3c99;
mem_array[45659] = 16'h4650;
mem_array[45658] = 16'hbd78;
mem_array[45661] = 16'h741b;
mem_array[45660] = 16'hbe2d;
mem_array[45663] = 16'hcb34;
mem_array[45662] = 16'h3f54;
mem_array[45665] = 16'h1296;
mem_array[45664] = 16'h3e22;
mem_array[45667] = 16'ha7e9;
mem_array[45666] = 16'hbb31;
mem_array[45669] = 16'hef70;
mem_array[45668] = 16'h3f4e;
mem_array[45671] = 16'h488e;
mem_array[45670] = 16'hbd59;
mem_array[45673] = 16'hb86b;
mem_array[45672] = 16'hbdda;
mem_array[45675] = 16'he6fc;
mem_array[45674] = 16'hbdc6;
mem_array[45677] = 16'hb1dd;
mem_array[45676] = 16'h3daa;
mem_array[45679] = 16'h2dda;
mem_array[45678] = 16'h3e3f;
mem_array[45681] = 16'h5d31;
mem_array[45680] = 16'h3db5;
mem_array[45683] = 16'hf450;
mem_array[45682] = 16'hbd98;
mem_array[45685] = 16'h0e7a;
mem_array[45684] = 16'hbd1c;
mem_array[45687] = 16'hfff5;
mem_array[45686] = 16'hbd2c;
mem_array[45689] = 16'h9a8b;
mem_array[45688] = 16'h3e92;
mem_array[45691] = 16'h127e;
mem_array[45690] = 16'hbf20;
mem_array[45693] = 16'h8d2f;
mem_array[45692] = 16'h3cf0;
mem_array[45695] = 16'hbcfd;
mem_array[45694] = 16'hbc5a;
mem_array[45697] = 16'hb768;
mem_array[45696] = 16'h3f37;
mem_array[45699] = 16'h7c1a;
mem_array[45698] = 16'h3ee7;
mem_array[45701] = 16'h657f;
mem_array[45700] = 16'hbe23;
mem_array[45703] = 16'hc183;
mem_array[45702] = 16'hbefc;
mem_array[45705] = 16'hdd65;
mem_array[45704] = 16'hbda1;
mem_array[45707] = 16'h39a7;
mem_array[45706] = 16'hbf47;
mem_array[45709] = 16'h4f87;
mem_array[45708] = 16'h3c28;
mem_array[45711] = 16'h4b71;
mem_array[45710] = 16'h3f73;
mem_array[45713] = 16'h50e5;
mem_array[45712] = 16'hbebf;
mem_array[45715] = 16'h7d89;
mem_array[45714] = 16'h3e93;
mem_array[45717] = 16'he9bf;
mem_array[45716] = 16'hbd9d;
mem_array[45719] = 16'h3218;
mem_array[45718] = 16'hbe2a;
mem_array[45721] = 16'h95a4;
mem_array[45720] = 16'hbbec;
mem_array[45723] = 16'h0abf;
mem_array[45722] = 16'h3f1b;
mem_array[45725] = 16'h4614;
mem_array[45724] = 16'h3dbd;
mem_array[45727] = 16'h3645;
mem_array[45726] = 16'hbe7f;
mem_array[45729] = 16'hb75b;
mem_array[45728] = 16'h3ec2;
mem_array[45731] = 16'he927;
mem_array[45730] = 16'hbe00;
mem_array[45733] = 16'h4a87;
mem_array[45732] = 16'hbe85;
mem_array[45735] = 16'h1841;
mem_array[45734] = 16'h3ca7;
mem_array[45737] = 16'ha2b3;
mem_array[45736] = 16'h3d11;
mem_array[45739] = 16'hb222;
mem_array[45738] = 16'h3e0c;
mem_array[45741] = 16'h8fa5;
mem_array[45740] = 16'hbda6;
mem_array[45743] = 16'h3b75;
mem_array[45742] = 16'h3dc8;
mem_array[45745] = 16'h41bf;
mem_array[45744] = 16'hbc4d;
mem_array[45747] = 16'hcd53;
mem_array[45746] = 16'hbd99;
mem_array[45749] = 16'h7e00;
mem_array[45748] = 16'h3e89;
mem_array[45751] = 16'h935b;
mem_array[45750] = 16'hbebf;
mem_array[45753] = 16'hc336;
mem_array[45752] = 16'hbd33;
mem_array[45755] = 16'h5765;
mem_array[45754] = 16'hbec0;
mem_array[45757] = 16'h9c11;
mem_array[45756] = 16'h3e20;
mem_array[45759] = 16'hd7e2;
mem_array[45758] = 16'h3dda;
mem_array[45761] = 16'h1326;
mem_array[45760] = 16'hbfac;
mem_array[45763] = 16'h2ea2;
mem_array[45762] = 16'h3dd1;
mem_array[45765] = 16'h7eb4;
mem_array[45764] = 16'h3c4f;
mem_array[45767] = 16'hfebe;
mem_array[45766] = 16'hbe8c;
mem_array[45769] = 16'hdc0c;
mem_array[45768] = 16'hbdb3;
mem_array[45771] = 16'h3fb6;
mem_array[45770] = 16'h3f0b;
mem_array[45773] = 16'h9dea;
mem_array[45772] = 16'h3d17;
mem_array[45775] = 16'h83f4;
mem_array[45774] = 16'h3def;
mem_array[45777] = 16'h5843;
mem_array[45776] = 16'h3c1e;
mem_array[45779] = 16'hbb23;
mem_array[45778] = 16'hbf1c;
mem_array[45781] = 16'h9075;
mem_array[45780] = 16'hbcb8;
mem_array[45783] = 16'h4912;
mem_array[45782] = 16'h3f1b;
mem_array[45785] = 16'h9ff8;
mem_array[45784] = 16'h3e37;
mem_array[45787] = 16'hb1da;
mem_array[45786] = 16'hbe11;
mem_array[45789] = 16'h018c;
mem_array[45788] = 16'h3e4c;
mem_array[45791] = 16'h7de3;
mem_array[45790] = 16'hbd8b;
mem_array[45793] = 16'hde16;
mem_array[45792] = 16'hbee3;
mem_array[45795] = 16'h22f6;
mem_array[45794] = 16'hbc26;
mem_array[45797] = 16'hbbfd;
mem_array[45796] = 16'hbd5f;
mem_array[45799] = 16'h6a7d;
mem_array[45798] = 16'h3de0;
mem_array[45801] = 16'h6d84;
mem_array[45800] = 16'hbcbf;
mem_array[45803] = 16'h5a96;
mem_array[45802] = 16'h3cc5;
mem_array[45805] = 16'h1b4f;
mem_array[45804] = 16'hbd8d;
mem_array[45807] = 16'hca1e;
mem_array[45806] = 16'hbd5e;
mem_array[45809] = 16'h9e2e;
mem_array[45808] = 16'h3e45;
mem_array[45811] = 16'h368b;
mem_array[45810] = 16'hbe80;
mem_array[45813] = 16'h1965;
mem_array[45812] = 16'h3d43;
mem_array[45815] = 16'h3d90;
mem_array[45814] = 16'hbed7;
mem_array[45817] = 16'h1282;
mem_array[45816] = 16'hbe0a;
mem_array[45819] = 16'hb1bc;
mem_array[45818] = 16'hbe20;
mem_array[45821] = 16'h40c0;
mem_array[45820] = 16'hbfb4;
mem_array[45823] = 16'h9a4f;
mem_array[45822] = 16'h3e46;
mem_array[45825] = 16'h197b;
mem_array[45824] = 16'h3d69;
mem_array[45827] = 16'h0f9e;
mem_array[45826] = 16'h3ead;
mem_array[45829] = 16'h2172;
mem_array[45828] = 16'hbd0c;
mem_array[45831] = 16'h9ed8;
mem_array[45830] = 16'h3e40;
mem_array[45833] = 16'h01d4;
mem_array[45832] = 16'h3e3f;
mem_array[45835] = 16'h1018;
mem_array[45834] = 16'h3e64;
mem_array[45837] = 16'hc843;
mem_array[45836] = 16'h3d99;
mem_array[45839] = 16'h2107;
mem_array[45838] = 16'hbf39;
mem_array[45841] = 16'h5ac8;
mem_array[45840] = 16'hbc55;
mem_array[45843] = 16'h99b2;
mem_array[45842] = 16'h3f2e;
mem_array[45845] = 16'h8299;
mem_array[45844] = 16'h3e62;
mem_array[45847] = 16'hb57e;
mem_array[45846] = 16'hbc11;
mem_array[45849] = 16'h62b0;
mem_array[45848] = 16'hbe19;
mem_array[45851] = 16'hf50a;
mem_array[45850] = 16'h3dba;
mem_array[45853] = 16'hb617;
mem_array[45852] = 16'hbed2;
mem_array[45855] = 16'h877c;
mem_array[45854] = 16'h3d7f;
mem_array[45857] = 16'h1dd4;
mem_array[45856] = 16'hbc8f;
mem_array[45859] = 16'hcf62;
mem_array[45858] = 16'h3ea3;
mem_array[45861] = 16'h2dff;
mem_array[45860] = 16'h3ce9;
mem_array[45863] = 16'hd61d;
mem_array[45862] = 16'h3c87;
mem_array[45865] = 16'h4bc9;
mem_array[45864] = 16'h3d26;
mem_array[45867] = 16'h54e2;
mem_array[45866] = 16'h3d16;
mem_array[45869] = 16'hd8c8;
mem_array[45868] = 16'hbd8c;
mem_array[45871] = 16'h5084;
mem_array[45870] = 16'hbec1;
mem_array[45873] = 16'h483d;
mem_array[45872] = 16'hbd18;
mem_array[45875] = 16'h2708;
mem_array[45874] = 16'hbee7;
mem_array[45877] = 16'hfd16;
mem_array[45876] = 16'h3d36;
mem_array[45879] = 16'h307d;
mem_array[45878] = 16'h3e3a;
mem_array[45881] = 16'hb2f9;
mem_array[45880] = 16'hbfb6;
mem_array[45883] = 16'he768;
mem_array[45882] = 16'h3de5;
mem_array[45885] = 16'hb4f3;
mem_array[45884] = 16'hbd90;
mem_array[45887] = 16'h2f31;
mem_array[45886] = 16'h3eba;
mem_array[45889] = 16'hd5a2;
mem_array[45888] = 16'hbca5;
mem_array[45891] = 16'h5151;
mem_array[45890] = 16'h3e0f;
mem_array[45893] = 16'h81e4;
mem_array[45892] = 16'h3e61;
mem_array[45895] = 16'h21ea;
mem_array[45894] = 16'h3e39;
mem_array[45897] = 16'h128d;
mem_array[45896] = 16'hbc66;
mem_array[45899] = 16'h94b3;
mem_array[45898] = 16'hbf59;
mem_array[45901] = 16'h295e;
mem_array[45900] = 16'h3f09;
mem_array[45903] = 16'h4eb2;
mem_array[45902] = 16'h3f78;
mem_array[45905] = 16'ha6c4;
mem_array[45904] = 16'h3f26;
mem_array[45907] = 16'h6fab;
mem_array[45906] = 16'hbe11;
mem_array[45909] = 16'hb612;
mem_array[45908] = 16'hbd99;
mem_array[45911] = 16'h106b;
mem_array[45910] = 16'hbcc4;
mem_array[45913] = 16'h393f;
mem_array[45912] = 16'h3d19;
mem_array[45915] = 16'h1edf;
mem_array[45914] = 16'h3eed;
mem_array[45917] = 16'he88c;
mem_array[45916] = 16'hbe2e;
mem_array[45919] = 16'hd4d9;
mem_array[45918] = 16'h3eac;
mem_array[45921] = 16'h0195;
mem_array[45920] = 16'h3c5b;
mem_array[45923] = 16'h3f15;
mem_array[45922] = 16'h3dd0;
mem_array[45925] = 16'h748f;
mem_array[45924] = 16'h3dae;
mem_array[45927] = 16'h5832;
mem_array[45926] = 16'hbdc8;
mem_array[45929] = 16'h8c3c;
mem_array[45928] = 16'hbe6a;
mem_array[45931] = 16'h17dd;
mem_array[45930] = 16'h3e52;
mem_array[45933] = 16'h819b;
mem_array[45932] = 16'hbab6;
mem_array[45935] = 16'h9589;
mem_array[45934] = 16'hbee7;
mem_array[45937] = 16'h45ff;
mem_array[45936] = 16'h3e63;
mem_array[45939] = 16'hac84;
mem_array[45938] = 16'h3e8d;
mem_array[45941] = 16'h9656;
mem_array[45940] = 16'hbfa6;
mem_array[45943] = 16'h2899;
mem_array[45942] = 16'hbf4a;
mem_array[45945] = 16'h15fe;
mem_array[45944] = 16'hbbb5;
mem_array[45947] = 16'h33a9;
mem_array[45946] = 16'hbd9d;
mem_array[45949] = 16'hf0a7;
mem_array[45948] = 16'hbdd3;
mem_array[45951] = 16'h5576;
mem_array[45950] = 16'h3e33;
mem_array[45953] = 16'h9e46;
mem_array[45952] = 16'hbe66;
mem_array[45955] = 16'h5b25;
mem_array[45954] = 16'hbe36;
mem_array[45957] = 16'hbaeb;
mem_array[45956] = 16'h3a44;
mem_array[45959] = 16'h37eb;
mem_array[45958] = 16'hbf5e;
mem_array[45961] = 16'h0c33;
mem_array[45960] = 16'h3e09;
mem_array[45963] = 16'h9a8e;
mem_array[45962] = 16'h3e16;
mem_array[45965] = 16'h3eda;
mem_array[45964] = 16'h3f43;
mem_array[45967] = 16'h09ed;
mem_array[45966] = 16'hbdd5;
mem_array[45969] = 16'h80ab;
mem_array[45968] = 16'h3f09;
mem_array[45971] = 16'haae1;
mem_array[45970] = 16'h3e83;
mem_array[45973] = 16'hdc22;
mem_array[45972] = 16'hbe0f;
mem_array[45975] = 16'h13ae;
mem_array[45974] = 16'h3f17;
mem_array[45977] = 16'hef51;
mem_array[45976] = 16'h3d66;
mem_array[45979] = 16'ha270;
mem_array[45978] = 16'h3e85;
mem_array[45981] = 16'h1334;
mem_array[45980] = 16'hbc60;
mem_array[45983] = 16'hcc97;
mem_array[45982] = 16'hbd18;
mem_array[45985] = 16'h3bc2;
mem_array[45984] = 16'h3dfc;
mem_array[45987] = 16'h61d9;
mem_array[45986] = 16'hbd31;
mem_array[45989] = 16'hcbd1;
mem_array[45988] = 16'hbe8e;
mem_array[45991] = 16'h8638;
mem_array[45990] = 16'h3e40;
mem_array[45993] = 16'hfadb;
mem_array[45992] = 16'h3c74;
mem_array[45995] = 16'hed68;
mem_array[45994] = 16'hbe76;
mem_array[45997] = 16'hf7e5;
mem_array[45996] = 16'h3ec3;
mem_array[45999] = 16'he393;
mem_array[45998] = 16'h3d8b;
mem_array[46001] = 16'h730f;
mem_array[46000] = 16'hbf61;
mem_array[46003] = 16'ha36f;
mem_array[46002] = 16'h3e42;
mem_array[46005] = 16'h8cf1;
mem_array[46004] = 16'h3d83;
mem_array[46007] = 16'hcb3b;
mem_array[46006] = 16'hbf4a;
mem_array[46009] = 16'h4c2a;
mem_array[46008] = 16'hbe78;
mem_array[46011] = 16'h7465;
mem_array[46010] = 16'h3f4b;
mem_array[46013] = 16'h7c72;
mem_array[46012] = 16'hbdf3;
mem_array[46015] = 16'ha239;
mem_array[46014] = 16'hbe70;
mem_array[46017] = 16'h5e3d;
mem_array[46016] = 16'hba82;
mem_array[46019] = 16'hd661;
mem_array[46018] = 16'hbf11;
mem_array[46021] = 16'hf9ec;
mem_array[46020] = 16'h3e07;
mem_array[46023] = 16'h2f9b;
mem_array[46022] = 16'hbe8f;
mem_array[46025] = 16'h06b4;
mem_array[46024] = 16'h3f5a;
mem_array[46027] = 16'h4bb3;
mem_array[46026] = 16'hbe04;
mem_array[46029] = 16'h0af3;
mem_array[46028] = 16'h3f43;
mem_array[46031] = 16'h45be;
mem_array[46030] = 16'h3e0a;
mem_array[46033] = 16'h6ac8;
mem_array[46032] = 16'hbecb;
mem_array[46035] = 16'ha024;
mem_array[46034] = 16'hbed2;
mem_array[46037] = 16'hd445;
mem_array[46036] = 16'hbf24;
mem_array[46039] = 16'h3aec;
mem_array[46038] = 16'h3e9b;
mem_array[46041] = 16'h5703;
mem_array[46040] = 16'hbdac;
mem_array[46043] = 16'h8c14;
mem_array[46042] = 16'h3c30;
mem_array[46045] = 16'h8274;
mem_array[46044] = 16'h3db2;
mem_array[46047] = 16'h89ef;
mem_array[46046] = 16'hbdf2;
mem_array[46049] = 16'h27bf;
mem_array[46048] = 16'hbee5;
mem_array[46051] = 16'hc181;
mem_array[46050] = 16'h3e83;
mem_array[46053] = 16'h2ff2;
mem_array[46052] = 16'hbd13;
mem_array[46055] = 16'h39cd;
mem_array[46054] = 16'hbed1;
mem_array[46057] = 16'hefe9;
mem_array[46056] = 16'h3c9d;
mem_array[46059] = 16'h564c;
mem_array[46058] = 16'hbe06;
mem_array[46061] = 16'hf2ba;
mem_array[46060] = 16'hbf7c;
mem_array[46063] = 16'h7b85;
mem_array[46062] = 16'h3e77;
mem_array[46065] = 16'hfeb0;
mem_array[46064] = 16'h3da4;
mem_array[46067] = 16'h365e;
mem_array[46066] = 16'h3e93;
mem_array[46069] = 16'h5ba7;
mem_array[46068] = 16'hbea9;
mem_array[46071] = 16'he483;
mem_array[46070] = 16'h3cbf;
mem_array[46073] = 16'he552;
mem_array[46072] = 16'h3cc9;
mem_array[46075] = 16'h6c8c;
mem_array[46074] = 16'hbe81;
mem_array[46077] = 16'hcf29;
mem_array[46076] = 16'hbdc1;
mem_array[46079] = 16'h5a18;
mem_array[46078] = 16'hbee4;
mem_array[46081] = 16'h9e52;
mem_array[46080] = 16'h3df1;
mem_array[46083] = 16'hf9b8;
mem_array[46082] = 16'h3f12;
mem_array[46085] = 16'h6bf6;
mem_array[46084] = 16'h3ee1;
mem_array[46087] = 16'hc213;
mem_array[46086] = 16'h3c40;
mem_array[46089] = 16'h8f37;
mem_array[46088] = 16'h3e31;
mem_array[46091] = 16'h7cd4;
mem_array[46090] = 16'h3e86;
mem_array[46093] = 16'hd6aa;
mem_array[46092] = 16'hbe81;
mem_array[46095] = 16'hd3d5;
mem_array[46094] = 16'hbd56;
mem_array[46097] = 16'h3263;
mem_array[46096] = 16'hbf13;
mem_array[46099] = 16'h9a94;
mem_array[46098] = 16'h3eca;
mem_array[46101] = 16'h2ecf;
mem_array[46100] = 16'hbd6f;
mem_array[46103] = 16'h4e83;
mem_array[46102] = 16'hbcd0;
mem_array[46105] = 16'h4d77;
mem_array[46104] = 16'h3e39;
mem_array[46107] = 16'hb8e3;
mem_array[46106] = 16'hbd88;
mem_array[46109] = 16'h2b5b;
mem_array[46108] = 16'hbe73;
mem_array[46111] = 16'h9b29;
mem_array[46110] = 16'hbeb7;
mem_array[46113] = 16'h23c8;
mem_array[46112] = 16'h3cc3;
mem_array[46115] = 16'hd80e;
mem_array[46114] = 16'hbec6;
mem_array[46117] = 16'h4fb5;
mem_array[46116] = 16'h3e92;
mem_array[46119] = 16'h2358;
mem_array[46118] = 16'h3f13;
mem_array[46121] = 16'h66b5;
mem_array[46120] = 16'hbf51;
mem_array[46123] = 16'h7420;
mem_array[46122] = 16'h3e01;
mem_array[46125] = 16'h5776;
mem_array[46124] = 16'h3cdb;
mem_array[46127] = 16'h2007;
mem_array[46126] = 16'h3b91;
mem_array[46129] = 16'h2b49;
mem_array[46128] = 16'hbea9;
mem_array[46131] = 16'h340e;
mem_array[46130] = 16'h3ef8;
mem_array[46133] = 16'hb276;
mem_array[46132] = 16'hbe1d;
mem_array[46135] = 16'hfd92;
mem_array[46134] = 16'hbdd0;
mem_array[46137] = 16'h57e7;
mem_array[46136] = 16'h3cc8;
mem_array[46139] = 16'hdd96;
mem_array[46138] = 16'hbf41;
mem_array[46141] = 16'h6315;
mem_array[46140] = 16'h3e9d;
mem_array[46143] = 16'ha25e;
mem_array[46142] = 16'h3ec8;
mem_array[46145] = 16'hcdc3;
mem_array[46144] = 16'h3eae;
mem_array[46147] = 16'hacae;
mem_array[46146] = 16'hbe1a;
mem_array[46149] = 16'he809;
mem_array[46148] = 16'h3ed8;
mem_array[46151] = 16'h3c6e;
mem_array[46150] = 16'h3e65;
mem_array[46153] = 16'hbdab;
mem_array[46152] = 16'hbde1;
mem_array[46155] = 16'h2cd8;
mem_array[46154] = 16'h3e64;
mem_array[46157] = 16'h65c1;
mem_array[46156] = 16'hbf28;
mem_array[46159] = 16'h9f58;
mem_array[46158] = 16'h3e53;
mem_array[46161] = 16'he42c;
mem_array[46160] = 16'h3bd0;
mem_array[46163] = 16'hd360;
mem_array[46162] = 16'h3b92;
mem_array[46165] = 16'h6109;
mem_array[46164] = 16'hbd5a;
mem_array[46167] = 16'h58d6;
mem_array[46166] = 16'hbb54;
mem_array[46169] = 16'ha2ab;
mem_array[46168] = 16'h3ce0;
mem_array[46171] = 16'he030;
mem_array[46170] = 16'hbeb6;
mem_array[46173] = 16'h8844;
mem_array[46172] = 16'hbe98;
mem_array[46175] = 16'ha5d0;
mem_array[46174] = 16'hbeec;
mem_array[46177] = 16'h5c40;
mem_array[46176] = 16'h3f28;
mem_array[46179] = 16'h3e36;
mem_array[46178] = 16'h3f81;
mem_array[46181] = 16'h326d;
mem_array[46180] = 16'hbfb6;
mem_array[46183] = 16'h64cc;
mem_array[46182] = 16'h3ec7;
mem_array[46185] = 16'h637c;
mem_array[46184] = 16'hbd83;
mem_array[46187] = 16'h0dfb;
mem_array[46186] = 16'hbdef;
mem_array[46189] = 16'h8694;
mem_array[46188] = 16'hbee8;
mem_array[46191] = 16'hc66e;
mem_array[46190] = 16'h3eaa;
mem_array[46193] = 16'h70d4;
mem_array[46192] = 16'hbcee;
mem_array[46195] = 16'h6567;
mem_array[46194] = 16'h3d35;
mem_array[46197] = 16'hd66e;
mem_array[46196] = 16'hbc51;
mem_array[46199] = 16'h568d;
mem_array[46198] = 16'hbf71;
mem_array[46201] = 16'h75a6;
mem_array[46200] = 16'h3f27;
mem_array[46203] = 16'hea78;
mem_array[46202] = 16'h3ed0;
mem_array[46205] = 16'ha22b;
mem_array[46204] = 16'h3e4f;
mem_array[46207] = 16'hd649;
mem_array[46206] = 16'hbea2;
mem_array[46209] = 16'h5711;
mem_array[46208] = 16'hbd88;
mem_array[46211] = 16'haf55;
mem_array[46210] = 16'h3e1c;
mem_array[46213] = 16'h1adf;
mem_array[46212] = 16'hbee6;
mem_array[46215] = 16'h6352;
mem_array[46214] = 16'hbed6;
mem_array[46217] = 16'hdf28;
mem_array[46216] = 16'hbef8;
mem_array[46219] = 16'he6e0;
mem_array[46218] = 16'h3e85;
mem_array[46221] = 16'ha3e0;
mem_array[46220] = 16'hbd32;
mem_array[46223] = 16'hcbea;
mem_array[46222] = 16'h3bae;
mem_array[46225] = 16'h1da4;
mem_array[46224] = 16'hbe2e;
mem_array[46227] = 16'hb3a7;
mem_array[46226] = 16'hbc98;
mem_array[46229] = 16'h4ea7;
mem_array[46228] = 16'hbea2;
mem_array[46231] = 16'hf134;
mem_array[46230] = 16'hbd10;
mem_array[46233] = 16'he99f;
mem_array[46232] = 16'hbe1b;
mem_array[46235] = 16'h065c;
mem_array[46234] = 16'hbf04;
mem_array[46237] = 16'hb5df;
mem_array[46236] = 16'h3f39;
mem_array[46239] = 16'hbe7f;
mem_array[46238] = 16'h3f86;
mem_array[46241] = 16'h34cc;
mem_array[46240] = 16'hc00c;
mem_array[46243] = 16'h9374;
mem_array[46242] = 16'h3f45;
mem_array[46245] = 16'h882a;
mem_array[46244] = 16'h3d81;
mem_array[46247] = 16'hb924;
mem_array[46246] = 16'hbe0b;
mem_array[46249] = 16'h150c;
mem_array[46248] = 16'hbeae;
mem_array[46251] = 16'h1506;
mem_array[46250] = 16'hbeb0;
mem_array[46253] = 16'h49ea;
mem_array[46252] = 16'h3ecd;
mem_array[46255] = 16'hc8de;
mem_array[46254] = 16'h3e04;
mem_array[46257] = 16'h6d86;
mem_array[46256] = 16'h3c82;
mem_array[46259] = 16'hcb6d;
mem_array[46258] = 16'hbfd9;
mem_array[46261] = 16'h0e14;
mem_array[46260] = 16'h3ddd;
mem_array[46263] = 16'h2e92;
mem_array[46262] = 16'hbe93;
mem_array[46265] = 16'he927;
mem_array[46264] = 16'h3d40;
mem_array[46267] = 16'hfaf4;
mem_array[46266] = 16'hbe71;
mem_array[46269] = 16'h49b0;
mem_array[46268] = 16'hbe67;
mem_array[46271] = 16'h63ea;
mem_array[46270] = 16'h3f3b;
mem_array[46273] = 16'h030b;
mem_array[46272] = 16'hbe62;
mem_array[46275] = 16'h68d1;
mem_array[46274] = 16'hbf52;
mem_array[46277] = 16'h5b37;
mem_array[46276] = 16'hbee2;
mem_array[46279] = 16'h3fe4;
mem_array[46278] = 16'h3e17;
mem_array[46281] = 16'h1b1c;
mem_array[46280] = 16'h3c85;
mem_array[46283] = 16'hd1d1;
mem_array[46282] = 16'h3da6;
mem_array[46285] = 16'h358e;
mem_array[46284] = 16'hbe0c;
mem_array[46287] = 16'hda76;
mem_array[46286] = 16'h3ce7;
mem_array[46289] = 16'h3e92;
mem_array[46288] = 16'hbdac;
mem_array[46291] = 16'h9ac1;
mem_array[46290] = 16'h3f52;
mem_array[46293] = 16'h4af0;
mem_array[46292] = 16'hbd5e;
mem_array[46295] = 16'h5620;
mem_array[46294] = 16'hbd38;
mem_array[46297] = 16'h086c;
mem_array[46296] = 16'h3f2c;
mem_array[46299] = 16'hb734;
mem_array[46298] = 16'hbef3;
mem_array[46301] = 16'hb9bf;
mem_array[46300] = 16'hbe28;
mem_array[46303] = 16'h8af6;
mem_array[46302] = 16'h3ee6;
mem_array[46305] = 16'h48fe;
mem_array[46304] = 16'h3d86;
mem_array[46307] = 16'h7851;
mem_array[46306] = 16'hbd56;
mem_array[46309] = 16'h6089;
mem_array[46308] = 16'hbe8a;
mem_array[46311] = 16'hae08;
mem_array[46310] = 16'hbf2d;
mem_array[46313] = 16'hb8fb;
mem_array[46312] = 16'h3f61;
mem_array[46315] = 16'h3664;
mem_array[46314] = 16'hbe1f;
mem_array[46317] = 16'he2da;
mem_array[46316] = 16'hbd63;
mem_array[46319] = 16'h0e45;
mem_array[46318] = 16'hbf22;
mem_array[46321] = 16'h18dd;
mem_array[46320] = 16'h3bfc;
mem_array[46323] = 16'he5b7;
mem_array[46322] = 16'h3ed3;
mem_array[46325] = 16'h1249;
mem_array[46324] = 16'h3e0d;
mem_array[46327] = 16'hff76;
mem_array[46326] = 16'hbe5f;
mem_array[46329] = 16'h5b10;
mem_array[46328] = 16'h3dae;
mem_array[46331] = 16'hb84e;
mem_array[46330] = 16'hbe4b;
mem_array[46333] = 16'h9bab;
mem_array[46332] = 16'h3d7c;
mem_array[46335] = 16'h4c82;
mem_array[46334] = 16'h3e14;
mem_array[46337] = 16'hbdb9;
mem_array[46336] = 16'hbe28;
mem_array[46339] = 16'hc994;
mem_array[46338] = 16'h3e99;
mem_array[46341] = 16'h0e77;
mem_array[46340] = 16'hbc8a;
mem_array[46343] = 16'hcfe6;
mem_array[46342] = 16'hbd93;
mem_array[46345] = 16'hfea6;
mem_array[46344] = 16'hbdd1;
mem_array[46347] = 16'h927b;
mem_array[46346] = 16'h3d00;
mem_array[46349] = 16'hf84e;
mem_array[46348] = 16'h3e41;
mem_array[46351] = 16'h5125;
mem_array[46350] = 16'h3f1e;
mem_array[46353] = 16'hf3d1;
mem_array[46352] = 16'hbc34;
mem_array[46355] = 16'hc930;
mem_array[46354] = 16'hbf10;
mem_array[46357] = 16'hcdb6;
mem_array[46356] = 16'h3e79;
mem_array[46359] = 16'h7136;
mem_array[46358] = 16'h3f22;
mem_array[46361] = 16'hd4c1;
mem_array[46360] = 16'hbf05;
mem_array[46363] = 16'he9fc;
mem_array[46362] = 16'hbd96;
mem_array[46365] = 16'h2e34;
mem_array[46364] = 16'hbda4;
mem_array[46367] = 16'h255d;
mem_array[46366] = 16'hbdb5;
mem_array[46369] = 16'h92d8;
mem_array[46368] = 16'h3e1d;
mem_array[46371] = 16'h0003;
mem_array[46370] = 16'h3f50;
mem_array[46373] = 16'h9622;
mem_array[46372] = 16'hbeea;
mem_array[46375] = 16'h2446;
mem_array[46374] = 16'hbdaf;
mem_array[46377] = 16'h4465;
mem_array[46376] = 16'h3b45;
mem_array[46379] = 16'hb67a;
mem_array[46378] = 16'hbdd5;
mem_array[46381] = 16'h6677;
mem_array[46380] = 16'h3e3a;
mem_array[46383] = 16'hfa3c;
mem_array[46382] = 16'h3ef5;
mem_array[46385] = 16'h4137;
mem_array[46384] = 16'hbe1d;
mem_array[46387] = 16'h5cb9;
mem_array[46386] = 16'h3e95;
mem_array[46389] = 16'hed4d;
mem_array[46388] = 16'hbe48;
mem_array[46391] = 16'hd7ae;
mem_array[46390] = 16'h3dfc;
mem_array[46393] = 16'h8c3d;
mem_array[46392] = 16'hbe7f;
mem_array[46395] = 16'he8c8;
mem_array[46394] = 16'hbe3d;
mem_array[46397] = 16'h5889;
mem_array[46396] = 16'hbeea;
mem_array[46399] = 16'hfda2;
mem_array[46398] = 16'h3ea6;
mem_array[46401] = 16'hb7bc;
mem_array[46400] = 16'hbcb8;
mem_array[46403] = 16'hd1df;
mem_array[46402] = 16'h3cce;
mem_array[46405] = 16'h2a50;
mem_array[46404] = 16'hbe0b;
mem_array[46407] = 16'h0006;
mem_array[46406] = 16'h3b85;
mem_array[46409] = 16'h7948;
mem_array[46408] = 16'h3f05;
mem_array[46411] = 16'h70cf;
mem_array[46410] = 16'h3e40;
mem_array[46413] = 16'he065;
mem_array[46412] = 16'hbe13;
mem_array[46415] = 16'h78cf;
mem_array[46414] = 16'hbf04;
mem_array[46417] = 16'hc35c;
mem_array[46416] = 16'h3f83;
mem_array[46419] = 16'h05dc;
mem_array[46418] = 16'h3e9e;
mem_array[46421] = 16'hdd85;
mem_array[46420] = 16'hbe3c;
mem_array[46423] = 16'h38b8;
mem_array[46422] = 16'hbebc;
mem_array[46425] = 16'he0ef;
mem_array[46424] = 16'h3d4c;
mem_array[46427] = 16'h83c9;
mem_array[46426] = 16'hbea9;
mem_array[46429] = 16'hbb76;
mem_array[46428] = 16'hbe5d;
mem_array[46431] = 16'ha89a;
mem_array[46430] = 16'h3ea6;
mem_array[46433] = 16'h5b6a;
mem_array[46432] = 16'hbe51;
mem_array[46435] = 16'h0cae;
mem_array[46434] = 16'hbef5;
mem_array[46437] = 16'ha052;
mem_array[46436] = 16'h3ddb;
mem_array[46439] = 16'h109f;
mem_array[46438] = 16'hbf6e;
mem_array[46441] = 16'he5e3;
mem_array[46440] = 16'h3e88;
mem_array[46443] = 16'hd934;
mem_array[46442] = 16'h3f7d;
mem_array[46445] = 16'hc662;
mem_array[46444] = 16'h3d11;
mem_array[46447] = 16'h2654;
mem_array[46446] = 16'h3eb5;
mem_array[46449] = 16'h57de;
mem_array[46448] = 16'hbe6d;
mem_array[46451] = 16'hd9b8;
mem_array[46450] = 16'hbca6;
mem_array[46453] = 16'hf757;
mem_array[46452] = 16'hbead;
mem_array[46455] = 16'h855f;
mem_array[46454] = 16'hbe67;
mem_array[46457] = 16'h6dc9;
mem_array[46456] = 16'hbe79;
mem_array[46459] = 16'h7c93;
mem_array[46458] = 16'hbe4a;
mem_array[46461] = 16'hc625;
mem_array[46460] = 16'hbdb8;
mem_array[46463] = 16'ha857;
mem_array[46462] = 16'hbd13;
mem_array[46465] = 16'hcb45;
mem_array[46464] = 16'hbe4b;
mem_array[46467] = 16'h69ed;
mem_array[46466] = 16'hbca0;
mem_array[46469] = 16'h6dce;
mem_array[46468] = 16'hbe29;
mem_array[46471] = 16'ha557;
mem_array[46470] = 16'hbe41;
mem_array[46473] = 16'hb8b7;
mem_array[46472] = 16'h3c83;
mem_array[46475] = 16'hda0b;
mem_array[46474] = 16'hbe93;
mem_array[46477] = 16'h748d;
mem_array[46476] = 16'h3f8f;
mem_array[46479] = 16'h156c;
mem_array[46478] = 16'hbdf8;
mem_array[46481] = 16'h52ee;
mem_array[46480] = 16'hbe85;
mem_array[46483] = 16'h5977;
mem_array[46482] = 16'h3cb0;
mem_array[46485] = 16'hd78f;
mem_array[46484] = 16'h3d0e;
mem_array[46487] = 16'h4569;
mem_array[46486] = 16'h3e97;
mem_array[46489] = 16'hd3d0;
mem_array[46488] = 16'h3e34;
mem_array[46491] = 16'h5150;
mem_array[46490] = 16'h3d08;
mem_array[46493] = 16'h182e;
mem_array[46492] = 16'hbea8;
mem_array[46495] = 16'h3b29;
mem_array[46494] = 16'hbf38;
mem_array[46497] = 16'hcfaa;
mem_array[46496] = 16'h3d59;
mem_array[46499] = 16'h191e;
mem_array[46498] = 16'hbf6c;
mem_array[46501] = 16'hb2e9;
mem_array[46500] = 16'h3e64;
mem_array[46503] = 16'h431b;
mem_array[46502] = 16'h3f00;
mem_array[46505] = 16'h8123;
mem_array[46504] = 16'h3cf2;
mem_array[46507] = 16'hb22e;
mem_array[46506] = 16'h3eac;
mem_array[46509] = 16'hb60c;
mem_array[46508] = 16'hbe58;
mem_array[46511] = 16'hd05a;
mem_array[46510] = 16'h3cc4;
mem_array[46513] = 16'hf747;
mem_array[46512] = 16'hbbed;
mem_array[46515] = 16'hf220;
mem_array[46514] = 16'hbd24;
mem_array[46517] = 16'h11fe;
mem_array[46516] = 16'hbdf7;
mem_array[46519] = 16'ha496;
mem_array[46518] = 16'h3e0c;
mem_array[46521] = 16'hf3c8;
mem_array[46520] = 16'hbc12;
mem_array[46523] = 16'h81b3;
mem_array[46522] = 16'h3c31;
mem_array[46525] = 16'h364f;
mem_array[46524] = 16'hbe07;
mem_array[46527] = 16'h11bf;
mem_array[46526] = 16'hbb06;
mem_array[46529] = 16'hbefa;
mem_array[46528] = 16'h3bdc;
mem_array[46531] = 16'ha9b0;
mem_array[46530] = 16'hbe45;
mem_array[46533] = 16'h8564;
mem_array[46532] = 16'hbde6;
mem_array[46535] = 16'hc65a;
mem_array[46534] = 16'hbecd;
mem_array[46537] = 16'h842f;
mem_array[46536] = 16'h3db5;
mem_array[46539] = 16'hbf63;
mem_array[46538] = 16'hbe40;
mem_array[46541] = 16'h022f;
mem_array[46540] = 16'hbf43;
mem_array[46543] = 16'ha87f;
mem_array[46542] = 16'hbdea;
mem_array[46545] = 16'h9aad;
mem_array[46544] = 16'h3d73;
mem_array[46547] = 16'h93af;
mem_array[46546] = 16'h3ed8;
mem_array[46549] = 16'hc62b;
mem_array[46548] = 16'hbf3b;
mem_array[46551] = 16'h903f;
mem_array[46550] = 16'hbcc1;
mem_array[46553] = 16'h7531;
mem_array[46552] = 16'h3ea8;
mem_array[46555] = 16'hbdd2;
mem_array[46554] = 16'h3eca;
mem_array[46557] = 16'h1bff;
mem_array[46556] = 16'h3caf;
mem_array[46559] = 16'h7355;
mem_array[46558] = 16'hbedc;
mem_array[46561] = 16'he516;
mem_array[46560] = 16'hbd22;
mem_array[46563] = 16'h9a9e;
mem_array[46562] = 16'h3e21;
mem_array[46565] = 16'h158a;
mem_array[46564] = 16'h3d03;
mem_array[46567] = 16'hcf55;
mem_array[46566] = 16'h3e57;
mem_array[46569] = 16'h874d;
mem_array[46568] = 16'hbd72;
mem_array[46571] = 16'hb066;
mem_array[46570] = 16'h3d07;
mem_array[46573] = 16'h705f;
mem_array[46572] = 16'h3dfe;
mem_array[46575] = 16'h4cc2;
mem_array[46574] = 16'hbd91;
mem_array[46577] = 16'hde34;
mem_array[46576] = 16'hbe1e;
mem_array[46579] = 16'h215d;
mem_array[46578] = 16'hbdd3;
mem_array[46581] = 16'hfd80;
mem_array[46580] = 16'h3c29;
mem_array[46583] = 16'h0f76;
mem_array[46582] = 16'h3cbc;
mem_array[46585] = 16'h5ed6;
mem_array[46584] = 16'hbdf0;
mem_array[46587] = 16'h5a8a;
mem_array[46586] = 16'h3ce4;
mem_array[46589] = 16'h3c67;
mem_array[46588] = 16'hbe50;
mem_array[46591] = 16'hbf68;
mem_array[46590] = 16'hbcbd;
mem_array[46593] = 16'h9da3;
mem_array[46592] = 16'hbd1e;
mem_array[46595] = 16'h26b7;
mem_array[46594] = 16'hbebf;
mem_array[46597] = 16'h74a5;
mem_array[46596] = 16'h3d09;
mem_array[46599] = 16'h04ad;
mem_array[46598] = 16'hbe66;
mem_array[46601] = 16'h7761;
mem_array[46600] = 16'hbe14;
mem_array[46603] = 16'h7ac5;
mem_array[46602] = 16'hbeda;
mem_array[46605] = 16'h8595;
mem_array[46604] = 16'h3d9b;
mem_array[46607] = 16'he0ac;
mem_array[46606] = 16'h3edc;
mem_array[46609] = 16'h345d;
mem_array[46608] = 16'hbf35;
mem_array[46611] = 16'hd65d;
mem_array[46610] = 16'hbe1b;
mem_array[46613] = 16'h435d;
mem_array[46612] = 16'hbef8;
mem_array[46615] = 16'h7183;
mem_array[46614] = 16'hbda4;
mem_array[46617] = 16'h77dd;
mem_array[46616] = 16'hbba1;
mem_array[46619] = 16'h3c4c;
mem_array[46618] = 16'h3c1e;
mem_array[46621] = 16'h67b6;
mem_array[46620] = 16'hbd5b;
mem_array[46623] = 16'hbd6d;
mem_array[46622] = 16'h3f43;
mem_array[46625] = 16'hcc27;
mem_array[46624] = 16'hbe46;
mem_array[46627] = 16'hd53f;
mem_array[46626] = 16'h3e32;
mem_array[46629] = 16'h8d4f;
mem_array[46628] = 16'h3eab;
mem_array[46631] = 16'h0b63;
mem_array[46630] = 16'h3d5d;
mem_array[46633] = 16'hcf95;
mem_array[46632] = 16'h3d97;
mem_array[46635] = 16'hfb87;
mem_array[46634] = 16'h3eec;
mem_array[46637] = 16'h98d1;
mem_array[46636] = 16'hbe12;
mem_array[46639] = 16'h4171;
mem_array[46638] = 16'hbc73;
mem_array[46641] = 16'hbdc0;
mem_array[46640] = 16'h3db6;
mem_array[46643] = 16'hc21a;
mem_array[46642] = 16'h3d0d;
mem_array[46645] = 16'h28fa;
mem_array[46644] = 16'hbf3c;
mem_array[46647] = 16'h3c97;
mem_array[46646] = 16'hbc34;
mem_array[46649] = 16'h6ec3;
mem_array[46648] = 16'hbd4b;
mem_array[46651] = 16'h21cc;
mem_array[46650] = 16'hbed6;
mem_array[46653] = 16'hfaed;
mem_array[46652] = 16'h3de8;
mem_array[46655] = 16'hadd1;
mem_array[46654] = 16'hbf08;
mem_array[46657] = 16'h2698;
mem_array[46656] = 16'h3eab;
mem_array[46659] = 16'h5644;
mem_array[46658] = 16'hbd88;
mem_array[46661] = 16'h6490;
mem_array[46660] = 16'hbf80;
mem_array[46663] = 16'h2a2b;
mem_array[46662] = 16'hbf33;
mem_array[46665] = 16'h1fa0;
mem_array[46664] = 16'h3d46;
mem_array[46667] = 16'h6507;
mem_array[46666] = 16'hbdd0;
mem_array[46669] = 16'hc2ce;
mem_array[46668] = 16'hbec4;
mem_array[46671] = 16'h85db;
mem_array[46670] = 16'hbe97;
mem_array[46673] = 16'h7d1b;
mem_array[46672] = 16'hbf1c;
mem_array[46675] = 16'h6361;
mem_array[46674] = 16'h3ef0;
mem_array[46677] = 16'h2c73;
mem_array[46676] = 16'h3c10;
mem_array[46679] = 16'hdef2;
mem_array[46678] = 16'hbe8d;
mem_array[46681] = 16'h4fe4;
mem_array[46680] = 16'h3d5a;
mem_array[46683] = 16'h3965;
mem_array[46682] = 16'h3edc;
mem_array[46685] = 16'h7f4a;
mem_array[46684] = 16'hbe16;
mem_array[46687] = 16'h4f3c;
mem_array[46686] = 16'h3d5e;
mem_array[46689] = 16'h91f4;
mem_array[46688] = 16'hbcfb;
mem_array[46691] = 16'hc103;
mem_array[46690] = 16'hbd6f;
mem_array[46693] = 16'h6577;
mem_array[46692] = 16'h3c86;
mem_array[46695] = 16'h24a4;
mem_array[46694] = 16'hbd06;
mem_array[46697] = 16'h3e5a;
mem_array[46696] = 16'hbde7;
mem_array[46699] = 16'hcd4b;
mem_array[46698] = 16'hbc88;
mem_array[46701] = 16'h440c;
mem_array[46700] = 16'h3cf7;
mem_array[46703] = 16'hf13a;
mem_array[46702] = 16'hbde5;
mem_array[46705] = 16'ha2f7;
mem_array[46704] = 16'hbdaa;
mem_array[46707] = 16'hb456;
mem_array[46706] = 16'h3ca9;
mem_array[46709] = 16'h2465;
mem_array[46708] = 16'h3d22;
mem_array[46711] = 16'h1141;
mem_array[46710] = 16'h3e3c;
mem_array[46713] = 16'hf95e;
mem_array[46712] = 16'hbd25;
mem_array[46715] = 16'h0a9e;
mem_array[46714] = 16'h3e9e;
mem_array[46717] = 16'h2450;
mem_array[46716] = 16'h3e57;
mem_array[46719] = 16'h0a0c;
mem_array[46718] = 16'h3e10;
mem_array[46721] = 16'h08e9;
mem_array[46720] = 16'hbc37;
mem_array[46723] = 16'hbdfc;
mem_array[46722] = 16'hbdd5;
mem_array[46725] = 16'h9650;
mem_array[46724] = 16'hbc03;
mem_array[46727] = 16'hbc96;
mem_array[46726] = 16'hbe77;
mem_array[46729] = 16'h6a12;
mem_array[46728] = 16'hbeb9;
mem_array[46731] = 16'haa03;
mem_array[46730] = 16'hbe93;
mem_array[46733] = 16'h39d8;
mem_array[46732] = 16'hbdba;
mem_array[46735] = 16'h5ccc;
mem_array[46734] = 16'h3e2b;
mem_array[46737] = 16'hc99b;
mem_array[46736] = 16'hbca1;
mem_array[46739] = 16'h2555;
mem_array[46738] = 16'hbdbf;
mem_array[46741] = 16'h30a6;
mem_array[46740] = 16'h3c96;
mem_array[46743] = 16'h9d09;
mem_array[46742] = 16'h3f06;
mem_array[46745] = 16'hf654;
mem_array[46744] = 16'hbd46;
mem_array[46747] = 16'h8e68;
mem_array[46746] = 16'hbc60;
mem_array[46749] = 16'he25b;
mem_array[46748] = 16'h3ea4;
mem_array[46751] = 16'h02f9;
mem_array[46750] = 16'hbd73;
mem_array[46753] = 16'hc50c;
mem_array[46752] = 16'h3d62;
mem_array[46755] = 16'h01cd;
mem_array[46754] = 16'h3e4f;
mem_array[46757] = 16'h2d10;
mem_array[46756] = 16'h3a1d;
mem_array[46759] = 16'h5fce;
mem_array[46758] = 16'hbbe2;
mem_array[46761] = 16'h9c14;
mem_array[46760] = 16'hbdc3;
mem_array[46763] = 16'h488c;
mem_array[46762] = 16'hbd81;
mem_array[46765] = 16'h4cb0;
mem_array[46764] = 16'h3ccd;
mem_array[46767] = 16'hb855;
mem_array[46766] = 16'hbd77;
mem_array[46769] = 16'h8cf4;
mem_array[46768] = 16'hbcbe;
mem_array[46771] = 16'h15ab;
mem_array[46770] = 16'hbed2;
mem_array[46773] = 16'h9a87;
mem_array[46772] = 16'h3d65;
mem_array[46775] = 16'hc444;
mem_array[46774] = 16'hbd72;
mem_array[46777] = 16'h1bb7;
mem_array[46776] = 16'h3eb9;
mem_array[46779] = 16'h83ea;
mem_array[46778] = 16'h3e0f;
mem_array[46781] = 16'ha563;
mem_array[46780] = 16'hbd97;
mem_array[46783] = 16'hed19;
mem_array[46782] = 16'hbe0f;
mem_array[46785] = 16'hd9e0;
mem_array[46784] = 16'h3be7;
mem_array[46787] = 16'h60f8;
mem_array[46786] = 16'hbef1;
mem_array[46789] = 16'h95c1;
mem_array[46788] = 16'h3d6c;
mem_array[46791] = 16'hc6bb;
mem_array[46790] = 16'h3ec9;
mem_array[46793] = 16'h8d41;
mem_array[46792] = 16'hbd9d;
mem_array[46795] = 16'h45e7;
mem_array[46794] = 16'h3eee;
mem_array[46797] = 16'h2877;
mem_array[46796] = 16'hbc88;
mem_array[46799] = 16'h23db;
mem_array[46798] = 16'hbeca;
mem_array[46801] = 16'hd7a8;
mem_array[46800] = 16'hbd78;
mem_array[46803] = 16'h1bf7;
mem_array[46802] = 16'h3c64;
mem_array[46805] = 16'h7a12;
mem_array[46804] = 16'h3cc5;
mem_array[46807] = 16'ha478;
mem_array[46806] = 16'hbc68;
mem_array[46809] = 16'h9e74;
mem_array[46808] = 16'hbb94;
mem_array[46811] = 16'h232e;
mem_array[46810] = 16'h3dd4;
mem_array[46813] = 16'hab3a;
mem_array[46812] = 16'h3d51;
mem_array[46815] = 16'hbfe1;
mem_array[46814] = 16'hbc40;
mem_array[46817] = 16'hb8f1;
mem_array[46816] = 16'h3cbe;
mem_array[46819] = 16'h885f;
mem_array[46818] = 16'hbbf1;
mem_array[46821] = 16'h600a;
mem_array[46820] = 16'h3c2b;
mem_array[46823] = 16'h3779;
mem_array[46822] = 16'hbc0a;
mem_array[46825] = 16'h95b1;
mem_array[46824] = 16'hbd57;
mem_array[46827] = 16'h95e0;
mem_array[46826] = 16'hbdc0;
mem_array[46829] = 16'hff70;
mem_array[46828] = 16'h3d8b;
mem_array[46831] = 16'hc4fd;
mem_array[46830] = 16'hbd80;
mem_array[46833] = 16'h294e;
mem_array[46832] = 16'hbb77;
mem_array[46835] = 16'h5fb6;
mem_array[46834] = 16'hbd10;
mem_array[46837] = 16'he922;
mem_array[46836] = 16'hbcf3;
mem_array[46839] = 16'h8ba5;
mem_array[46838] = 16'hbd59;
mem_array[46841] = 16'h86af;
mem_array[46840] = 16'h3d8a;
mem_array[46843] = 16'h6503;
mem_array[46842] = 16'h3c59;
mem_array[46845] = 16'h83ef;
mem_array[46844] = 16'hbce8;
mem_array[46847] = 16'h6832;
mem_array[46846] = 16'h3d25;
mem_array[46849] = 16'h27d1;
mem_array[46848] = 16'h3dc4;
mem_array[46851] = 16'h5257;
mem_array[46850] = 16'h3dcc;
mem_array[46853] = 16'hf0aa;
mem_array[46852] = 16'hbd2f;
mem_array[46855] = 16'hd8ef;
mem_array[46854] = 16'h3bab;
mem_array[46857] = 16'hab58;
mem_array[46856] = 16'h3d26;
mem_array[46859] = 16'hcc07;
mem_array[46858] = 16'h3b79;
mem_array[46861] = 16'haa9a;
mem_array[46860] = 16'hbd2d;
mem_array[46863] = 16'hcbf2;
mem_array[46862] = 16'hbd56;
mem_array[46865] = 16'h0b43;
mem_array[46864] = 16'h3ddc;
mem_array[46867] = 16'h7ac9;
mem_array[46866] = 16'hbd39;
mem_array[46869] = 16'h01ae;
mem_array[46868] = 16'h3c06;
mem_array[46871] = 16'hb8e6;
mem_array[46870] = 16'hbcfa;
mem_array[46873] = 16'h8b68;
mem_array[46872] = 16'hbd86;
mem_array[46875] = 16'he5cd;
mem_array[46874] = 16'hbd8f;
mem_array[46877] = 16'h40f5;
mem_array[46876] = 16'h3bda;
mem_array[46879] = 16'ha362;
mem_array[46878] = 16'h3cf6;
mem_array[46881] = 16'h35bf;
mem_array[46880] = 16'h3d92;
mem_array[46883] = 16'hea15;
mem_array[46882] = 16'hbd1f;
mem_array[46885] = 16'h3005;
mem_array[46884] = 16'h3d16;
mem_array[46887] = 16'hc23a;
mem_array[46886] = 16'h3d1e;
mem_array[46889] = 16'hb342;
mem_array[46888] = 16'hbc5c;
mem_array[46891] = 16'h45c3;
mem_array[46890] = 16'h3961;
mem_array[46893] = 16'hf8da;
mem_array[46892] = 16'hbd00;
mem_array[46895] = 16'hb723;
mem_array[46894] = 16'hbd39;
mem_array[46897] = 16'hb638;
mem_array[46896] = 16'h3d1f;
mem_array[46899] = 16'h09fb;
mem_array[46898] = 16'hbd2f;
mem_array[46901] = 16'h6aa8;
mem_array[46900] = 16'hbde4;
mem_array[46903] = 16'h07bc;
mem_array[46902] = 16'hbbd1;
mem_array[46905] = 16'h1136;
mem_array[46904] = 16'hbb84;
mem_array[46907] = 16'h296e;
mem_array[46906] = 16'hbce9;
mem_array[46909] = 16'h1bee;
mem_array[46908] = 16'h3de6;
mem_array[46911] = 16'h1369;
mem_array[46910] = 16'hbd0b;
mem_array[46913] = 16'hc021;
mem_array[46912] = 16'h3db3;
mem_array[46915] = 16'h986d;
mem_array[46914] = 16'hbca0;
mem_array[46917] = 16'h50da;
mem_array[46916] = 16'h3d7d;
mem_array[46919] = 16'h8006;
mem_array[46918] = 16'hbd19;
mem_array[46921] = 16'hb674;
mem_array[46920] = 16'h3d93;
mem_array[46923] = 16'heac9;
mem_array[46922] = 16'hbaef;
mem_array[46925] = 16'hdcaa;
mem_array[46924] = 16'hbc5f;
mem_array[46927] = 16'he46d;
mem_array[46926] = 16'h3d31;
mem_array[46929] = 16'h0f6a;
mem_array[46928] = 16'hbd3c;
mem_array[46931] = 16'hcc60;
mem_array[46930] = 16'h3d0c;
mem_array[46933] = 16'hdfb6;
mem_array[46932] = 16'h3d9a;
mem_array[46935] = 16'h2b6c;
mem_array[46934] = 16'hbd31;
mem_array[46937] = 16'h20f4;
mem_array[46936] = 16'hbd71;
mem_array[46939] = 16'hae9b;
mem_array[46938] = 16'hbb42;
mem_array[46941] = 16'haea3;
mem_array[46940] = 16'h3d3d;
mem_array[46943] = 16'h0088;
mem_array[46942] = 16'h3dab;
mem_array[46945] = 16'h5aba;
mem_array[46944] = 16'hbd73;
mem_array[46947] = 16'h7f7c;
mem_array[46946] = 16'h3d66;
mem_array[46949] = 16'h9db5;
mem_array[46948] = 16'hbd65;
mem_array[46951] = 16'h2380;
mem_array[46950] = 16'hbd64;
mem_array[46953] = 16'h00dc;
mem_array[46952] = 16'h3c39;
mem_array[46955] = 16'he3d3;
mem_array[46954] = 16'h3c9d;
mem_array[46957] = 16'h5b31;
mem_array[46956] = 16'h3d94;
mem_array[46959] = 16'h2bd9;
mem_array[46958] = 16'hbbb2;
mem_array[46961] = 16'h30dd;
mem_array[46960] = 16'hbde8;
mem_array[46963] = 16'h498f;
mem_array[46962] = 16'h3cb4;
mem_array[46965] = 16'h81e0;
mem_array[46964] = 16'hbd93;
mem_array[46967] = 16'hbb4f;
mem_array[46966] = 16'hbd37;
mem_array[46969] = 16'h328f;
mem_array[46968] = 16'hbcab;
mem_array[46971] = 16'h31c2;
mem_array[46970] = 16'h3d64;
mem_array[46973] = 16'h6e47;
mem_array[46972] = 16'h3d1e;
mem_array[46975] = 16'h3806;
mem_array[46974] = 16'h3bf2;
mem_array[46977] = 16'hc236;
mem_array[46976] = 16'hbd84;
mem_array[46979] = 16'h543b;
mem_array[46978] = 16'h3d23;
mem_array[46981] = 16'h86e1;
mem_array[46980] = 16'hbd9c;
mem_array[46983] = 16'h6faf;
mem_array[46982] = 16'h3d7c;
mem_array[46985] = 16'h3baf;
mem_array[46984] = 16'h3b9f;
mem_array[46987] = 16'h0ebb;
mem_array[46986] = 16'hbd90;
mem_array[46989] = 16'h5598;
mem_array[46988] = 16'hba35;
mem_array[46991] = 16'hcb2f;
mem_array[46990] = 16'hbd43;
mem_array[46993] = 16'h3634;
mem_array[46992] = 16'hbcd1;
mem_array[46995] = 16'hc1e2;
mem_array[46994] = 16'hbd0f;
mem_array[46997] = 16'hf273;
mem_array[46996] = 16'h3dd9;
mem_array[46999] = 16'h5bc1;
mem_array[46998] = 16'hbdad;
mem_array[47001] = 16'h1ee8;
mem_array[47000] = 16'hbc3d;
mem_array[47003] = 16'hd747;
mem_array[47002] = 16'hbd01;
mem_array[47005] = 16'h3992;
mem_array[47004] = 16'h3d7c;
mem_array[47007] = 16'h514a;
mem_array[47006] = 16'hbc66;
mem_array[47009] = 16'he8d5;
mem_array[47008] = 16'hbd5c;
mem_array[47011] = 16'h6900;
mem_array[47010] = 16'h3cc7;
mem_array[47013] = 16'hfde7;
mem_array[47012] = 16'h3d49;
mem_array[47015] = 16'h966a;
mem_array[47014] = 16'hbd57;
mem_array[47017] = 16'h2830;
mem_array[47016] = 16'hbd20;
mem_array[47019] = 16'hce81;
mem_array[47018] = 16'hbd56;
mem_array[47021] = 16'ha16a;
mem_array[47020] = 16'h3ca0;
mem_array[47023] = 16'h40c4;
mem_array[47022] = 16'hbd4c;
mem_array[47025] = 16'hff73;
mem_array[47024] = 16'hbcf2;
mem_array[47027] = 16'hcb48;
mem_array[47026] = 16'hbc6b;
mem_array[47029] = 16'h2812;
mem_array[47028] = 16'hbdd5;
mem_array[47031] = 16'h2b10;
mem_array[47030] = 16'h3d46;
mem_array[47033] = 16'h2175;
mem_array[47032] = 16'hbc80;
mem_array[47035] = 16'hf18b;
mem_array[47034] = 16'h3dda;
mem_array[47037] = 16'h45a5;
mem_array[47036] = 16'hbd94;
mem_array[47039] = 16'h16d3;
mem_array[47038] = 16'hbdad;


endtask

endmodule