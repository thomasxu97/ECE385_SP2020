module weight_mat_w2(
	input [8:0] addr,
	output [31:0] weight
);
	parameter ADDR_WIDTH = 9;
   parameter DATA_WIDTH = 32;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	32'h3C25EF22,
32'hBDD77885,
32'hBE915F81,
32'h3EAD9289,
32'h3E020F09,
32'h3D651423,
32'h3A2A886,
32'h3F63C5E0,
32'h3EF90CF9,
32'hBDC0A10E,
32'h3F9746F7,
32'h3F27C8F4,
32'hBF5E6FDD,
32'h3FAAD3BE,
32'hBF03B8DF,
32'h3E5347B9,
32'hBF3289D9,
32'h3FD5D5A9,
32'h3F56B591,
32'h3EAB82F1,
32'h3F099D8B,
32'h3F152E9B,
32'h3F13AA9B,
32'hBEE8BEC2,
32'h3D25B162,
32'hBF792CC1,
32'hBD38B5CE,
32'h3F199DB3,
32'h3F412D50,
32'h3F2B2668,
32'h3E3EB84F,
32'h3F494F4A,
32'h3F10F951,
32'h3E843884,
32'hBD639966,
32'h3E070864,
32'hBCC4CAC3,
32'hBD070E39,
32'hBEB8A68F,
32'h3DFD5C9A,
32'hBF550B29,
32'hBE0B99D9,
32'h3F4910D6,
32'h3EB21DAC,
32'hBE5FC9C7,
32'h3CDB8E99,
32'h3DEAF2E5,
32'hBE9D019A,
32'h3F18D38C,
32'hBCAA31D4,
32'hBCDCD4BA,
32'hBE1ECF13,
32'hBF2FF789,
32'hBF2A70C1,
32'hBD1A4FB2,
32'hBE8C3838,
32'h3E10D04E,
32'hBE87EB25,
32'hBE3BDA14,
32'hBEF79252,
32'hBCDFEFE5,
32'hBEEE0E2B,
32'h3F49D8F0,
32'h3F029A1D,
32'h3D1E6DEE,
32'h3DD500F3,
32'h3D81C371,
32'h3E1825AA,
32'hBEE6B244,
32'hBEACE7A1,
32'h3F1D5CE9,
32'h3F00B63E,
32'h175F7BFE,
32'h3E94A637,
32'hBE079915,
32'h3C1255D9,
32'hBDDF35AC,
32'hBEE86B57,
32'h3EAFCD20,
32'hBCA96208,
32'hBF9BDB48,
32'h3DED68AA,
32'h3EE90C3F,
32'h3F1E778B,
32'hBDBFF698,
32'h3F164FD4,
32'hBC1A6075,
32'hBF2A2F1C,
32'h3F5A75C3,
32'hBE95CBDD,
32'h3D80C3A4,
32'h3DC384A9,
32'h3EC2F15A,
32'hBEFFADE7,
32'hBD22AB21,
32'h3C877BE6,
32'h3D30481C,
32'hBF11F5ED,
32'hBE6399A1,
32'h3DBAA969,
32'hBE95626D,
32'hBE98E75D,
32'h3EAE4D8F,
32'hBDDBDF0A,
32'h3F232DFA,
32'h3D28A5CE,
32'h3D8BB51E,
32'h3F23F6BD,
32'h3E91BA33,
32'hBDCD577B,
32'hBD26A415,
32'h3E673D3C,
32'hBEF7371D,
32'h3EC992CE,
32'h3D62A245,
32'hBE025CFC,
32'hBEF5ECCF,
32'hBE4AF8ED,
32'hBEA9718C,
32'h3F4242C9,
32'h3EA83224,
32'h3F8B37C8,
32'h3E9374CD,
32'h3E28E0AA,
32'h1DDD86E8,
32'h3E2014F8,
32'h3D11D38E,
32'h3ECB03F4,
32'h3DD8280F,
32'h3F244B61,
32'hBFC06298,
32'hBF36F1EC,
32'h3F994FB7,
32'h3E7E5008,
32'h3E8B7AE2,
32'h3D797DE2,
32'h3EB4CA4F,
32'hBF9B129F,
32'h3DCACA47,
32'h3E09171A,
32'h3D2FB713,
32'hBDC165A1,
32'h3F579006,
32'hBF3BA61C,
32'h3D009FA3,
32'h3F5E9585,
32'h3EB8C979,
32'hBE169C2B,
32'h3F9B5FCD,
32'hBF5DA521,
32'hBD7DAA61,
32'h3E69FC85,
32'h3F10508C,
32'h3E430602,
32'hBD3C8730,
32'h3E135366,
32'hBE4077C8,
32'hBEE30E12,
32'h3E7941CC,
32'hBF0B7E99,
32'h3D8DE9B2,
32'h3E63CAA3,
32'h3D166B4A,
32'hBEA7F2CC,
32'h3D01602C,
32'h3ED4D068,
32'h3E44463D,
32'hBCC78930,
32'h3C03F1D2,
32'hBD2AA3D4,
32'h3E64125E,
32'h3E636227,
32'h3D8EDB59,
32'hBD861B0B,
32'h3E2BB2E1,
32'h3E88274E,
32'hBE3F34BA,
32'hBEAC06C3,
32'h3CA1922C,
32'h0EDB9EB4,
32'hBC91C987,
32'h3E1D6E82,
32'hBF417E98,
32'h3E2775D4,
32'hBF001202,
32'hBDE4ABFB,
32'hBE4DFD38,
32'hBEAD31CB,
32'h3E87FB4B,
32'h1753ACDB,
32'hBCCF5D29,
32'hBE48A528,
32'h3ED99A76,
32'h3E4787C5,
32'hBEA0CA73,
32'h3E831F92,
32'h3F86334E,
32'hBE8165EC,
32'hBF6F23B5,
32'hBEB3EC64,
32'h3DD70926,
32'hBDC1231D,
32'h3E6DCAAF,
32'hBD867AA2,
32'h3F02D2C0,
32'hBE215605,
32'hBF16D7C9,
32'h3FBD9FEB,
32'h3F0186D9,
32'hBE05847A,
32'h3E355FFB,
32'h3F300C55,
32'h3E13B756,
32'hBEFD513C,
32'hBD50F309,
32'h3E070BE4,
32'h3D029504,
32'h3EB91593,
32'hBD5FCBC2,
32'h3EB50B59,
32'hBE843978,
32'hBE9BB95D,
32'h3F23E27B,
32'h3F446265,
32'h3E573279,
32'h1DD93DCE,
32'hBE76B85E,
32'hBEB78506,
32'hBE02F594,
32'h3D01FBB5,
32'h5DE44793,
32'hBD3F8D7F,
32'h3E356461,
32'hBF4278AE,
32'h3D299C50,
32'hBEC37052,
32'hBD1345C2,
32'hBD5A1347,
32'hBE4FC568,
32'hBCE9B764,
32'h3E7AED23,
32'h3F750661,
32'hBF556F4A,
32'hBEFFE5DF,
32'hBE05FDB2,
32'hBDD41F8D,
32'hBD4904F8,
32'h3E69300E,
32'hBF6C41FE,
32'h3F046A33,
32'h3EB415FB,
32'hBE0BF9D4,
32'h3F07A9BC,
32'h3F200D23,
32'hBE4B4070,
32'hBD1F8815,
32'h3D0ED2B8,
32'hBFB36087,
32'hBF8B5A68,
32'hBE863179,
32'h3E263DFE,
32'hBE9F186E,
32'hBF2ABF2B,
32'hBE990511,
32'hBE9E313F,
32'h3E292A35,
32'h3F5D131D,
32'h3EC72F93,
32'h3F1CE7E4,
32'hBF0816E0,
32'hBD1781AE,
32'hBEEC59EC,
32'h3F28F843,
32'h3EB26F74,
32'h3DABD011,
32'h3D4089FE,
32'h3DA31C3D,
32'hBE460596,
32'hBEA36724,
32'hBE96F2FF,
32'h3ECFD208,
32'h3E4F47EA,
32'hBE4397C0,
32'hBDA044E6,
32'hBECB1A1B,
32'hBD91E7B0,
32'hBEE7F5CA,
32'hBE1F8214,
32'hBEF5AC95,
32'h3CB6BB98,
32'h3E373DE3,
32'hBC4152D1,
32'hBE8CDCB2,
32'h3EC15DE2,
32'hBED2E6C1,
32'h3F125979,
32'h3F2F246B,
32'h3E1815D6,
32'h3E8E3889,
32'h3E778577,
32'hBD757CFD,
32'hBD84DEF5,
32'hBF502920,
32'hBF2DBB38,
32'hBE183986,
32'h3E273252,
32'hBDE55AD8,
32'hBF50FE47,
32'hBEEA3C34,
32'hBEED5CF9,
32'h3ECB130F,
32'h3F1FE341,
32'h3EF8CE9D,
32'h3E6A844C,
32'hBF14BE5B,
32'h1DE625A4,
32'hBEAD114E,
32'hBF240CFD,
32'hBE9A31A0,
32'h2ED77A1A,
32'h075821C7,
32'h3CAC33BE,
32'hBEEBA4F2,
32'hBD521BC8,
32'hBC95E25C,
32'hBF09C0E0,
32'hBE427766,
32'hBF4C75DA,
32'hBF2D6905,
32'hBE918BFC,
32'hBEEAA14C,
32'hBF227B57,
32'h3F181BE6,
32'h3E9875BE,
32'hBF846EE8,
32'hBF242B96,
32'hBE95567F,
32'hBFCA8A10,
32'h3EC1A6FB,
32'hBF8C54C8,
32'hBF5B7B38,
32'hBED4B519,
32'h3F396E5B,
32'hBF448FCE,
32'hBF67BAA7,
32'hBC5CDF91,
32'hBD59A359,
32'hBDB1F1A4,
32'hBDCF8C51,
32'hBD32C7A4,
32'hBCA8AD50,
32'h5DF59330,
32'hBE7DF495,
32'hBF03A693,
32'hBDAD9564,
32'hBE90181D,
32'hBE6FCA06,
32'h3D7D90F6,
32'hBEDF886C,
32'hBF13F17F,
32'h3DC4DED0,
32'h3E6EC3A0,
32'h3F135A42,
32'h3E0E63F4,
32'hBD170A0A,
32'h3D056092,
32'h3E00B9D2,
32'hBEA19ECE,
32'h3DC2F084,
32'h3DB9670C,
32'hBF42D175,
32'hBE2BF50B,
32'h3E8A1FD4,
32'hBD2E4173,
32'h3F428526,
32'h3E2E0023,
32'hBED58F47,
32'h3F7A734C,
32'h3F31F941,
32'h3E245EE8,
32'h3ED0F118,
32'h3EB6C98E,
32'h3EE2CDB9,
32'hBEF61837,
32'hBDD6EB34,
32'hBF15A645,
32'h3D78C4AF,
32'h3EC5A213,
32'h3ECB6BB6,
32'h3E963B8B,
32'h1755ECB6,
32'hBDC05069,
32'hBEBEF5B9,
32'hBE68DB09,
32'h5DC0C38D,
32'hBD55D4A4,
32'h3A4A42A,
32'hBE3FB262,
32'h3E81F9EC,
32'h3CBE3EC1,
32'hBE1EA538,
32'hBF10371B,
32'hBE3E6AE4,
32'hBF01E152,
32'h3D8ECBB1,
32'h3A2C2EE,
32'hBDABA94A,
32'hBE99ADDE,
32'hBE8280DD,
32'hBDC33526,
32'hBF998C0A,
32'h3E64AFCD,
32'hBF9F2282,
32'h3F91AA3A,
32'hBDE78FCE,
32'h3E5AD414,
32'hBFD788D8,
32'hBE90675C,
32'h3C3CA1E7,
32'h3D3A9627,
32'h3E5ACB4D,
32'h3F313667,
32'hBE59CA3F,
32'hBE0CCF34,
32'hBF413DEA,
32'hBD417091,
32'hBC910AF4,
32'h3E901EC0,
32'hBEDCE184,
32'h3F36D265,
32'h3E886197,
32'hBF2F7999,
32'h3F9658D8,
32'h3F19F43F,
32'h3EF233B6,
32'hBD058E57,
32'h3C8AB14D,
32'hBE83CC8E,
32'hBF0985BF,
32'hBDD60CFA,
32'h3CDEA670,
32'hBE05A1B8,
32'hBE4A4A40,
32'hBE588FEE,
32'hBD9349CE,
32'hBF4AFF83,
32'h3E3C8059,
32'hBF02D1F9,
32'hBEB7417B,
32'hBE8AF785
};
	assign weight = ROM[addr];
endmodule
