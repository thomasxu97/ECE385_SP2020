module font_rom ( input [10:0]	addr,
						output [7:0]	data
					 );

	parameter ADDR_WIDTH = 11;
   parameter DATA_WIDTH =  8;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x01
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111110, // 2  ******
        8'b10000001, // 3 *      *
        8'b10100101, // 4 * *  * *
        8'b10000001, // 5 *      *
        8'b10000001, // 6 *      *
        8'b10111101, // 7 * **** *
        8'b10011001, // 8 *  **  *
        8'b10000001, // 9 *      *
        8'b10000001, // a *      *
        8'b01111110, // b  ******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x02
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111110, // 2  ******
        8'b11111111, // 3 ********
        8'b11011011, // 4 ** ** **
        8'b11111111, // 5 ********
        8'b11111111, // 6 ********
        8'b11000011, // 7 **    **
        8'b11100111, // 8 ***  ***
        8'b11111111, // 9 ********
        8'b11111111, // a ********
        8'b01111110, // b  ******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x03
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00110110, // 4  ** **
        8'b01111111, // 5 *******
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01111111, // 8 *******
        8'b00111110, // 9  *****
        8'b00011100, // a   ***
        8'b00001000, // b    *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x04
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00001000, // 4    *
        8'b00011100, // 5   ***
        8'b00111110, // 6  *****
        8'b01111111, // 7 *******
        8'b00111110, // 8  *****
        8'b00011100, // 9   ***
        8'b00001000, // a    *
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x05
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00011000, // 3    **
        8'b00111100, // 4   ****
        8'b00111100, // 5   ****
        8'b11100111, // 6 ***  ***
        8'b11100111, // 7 ***  ***
        8'b11100111, // 8 ***  ***
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x06
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00011000, // 3    **
        8'b00111100, // 4   ****
        8'b01111110, // 5  ******
        8'b11111111, // 6 ********
        8'b11111111, // 7 ********
        8'b01111110, // 8  ******
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x07
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00011000, // 6    **
        8'b00111100, // 7   ****
        8'b00111100, // 8   ****
        8'b00011000, // 9    **
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x08
        8'b11111111, // 0 ********
        8'b11111111, // 1 ********
        8'b11111111, // 2 ********
        8'b11111111, // 3 ********
        8'b11111111, // 4 ********
        8'b11111111, // 5 ********
        8'b11100111, // 6 ***  ***
        8'b11000011, // 7 **    **
        8'b11000011, // 8 **    **
        8'b11100111, // 9 ***  ***
        8'b11111111, // a ********
        8'b11111111, // b ********
        8'b11111111, // c ********
        8'b11111111, // d ********
        8'b11111111, // e ********
        8'b11111111, // f ********
         // code x09
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111100, // 5   ****
        8'b01100110, // 6  **  **
        8'b01000010, // 7  *    *
        8'b01000010, // 8  *    *
        8'b01100110, // 9  **  **
        8'b00111100, // a   ****
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x0a
        8'b11111111, // 0 ********
        8'b11111111, // 1 ********
        8'b11111111, // 2 ********
        8'b11111111, // 3 ********
        8'b11111111, // 4 ********
        8'b11000011, // 5 **    **
        8'b10011001, // 6 *  **  *
        8'b10111101, // 7 * **** *
        8'b10111101, // 8 * **** *
        8'b10011001, // 9 *  **  *
        8'b11000011, // a **    **
        8'b11111111, // b ********
        8'b11111111, // c ********
        8'b11111111, // d ********
        8'b11111111, // e ********
        8'b11111111, // f ********
         // code x0b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111000, // 2    ****
        8'b01110000, // 3     ***
        8'b01011000, // 4    ** *
        8'b01001100, // 5   **  *
        8'b00011110, // 6  ****
        8'b00110011, // 7 **  **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b00011110, // b  ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x0c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b01100110, // 6  **  **
        8'b00111100, // 7   ****
        8'b00011000, // 8    **
        8'b01111110, // 9  ******
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x0d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111100, // 2   ******
        8'b11001100, // 3   **  **
        8'b11111100, // 4   ******
        8'b00001100, // 5   **
        8'b00001100, // 6   **
        8'b00001100, // 7   **
        8'b00001100, // 8   **
        8'b00001110, // 9  ***
        8'b00001111, // a ****
        8'b00000111, // b ***
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x0e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2  *******
        8'b11000110, // 3  **   **
        8'b11111110, // 4  *******
        8'b11000110, // 5  **   **
        8'b11000110, // 6  **   **
        8'b11000110, // 7  **   **
        8'b11000110, // 8  **   **
        8'b11100110, // 9  **  ***
        8'b11100111, // a ***  ***
        8'b01100111, // b ***  **
        8'b00000011, // c **
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x0f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b11011011, // 5 ** ** **
        8'b00111100, // 6   ****
        8'b11100111, // 7 ***  ***
        8'b00111100, // 8   ****
        8'b11011011, // 9 ** ** **
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x10
        8'b00000000, // 0
        8'b00000001, // 1 *
        8'b00000011, // 2 **
        8'b00000111, // 3 ***
        8'b00001111, // 4 ****
        8'b00011111, // 5 *****
        8'b01111111, // 6 *******
        8'b00011111, // 7 *****
        8'b00001111, // 8 ****
        8'b00000111, // 9 ***
        8'b00000011, // a **
        8'b00000001, // b *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x11
        8'b00000000, // 0
        8'b01000000, // 1       *
        8'b01100000, // 2      **
        8'b01110000, // 3     ***
        8'b01111000, // 4    ****
        8'b01111100, // 5   *****
        8'b01111111, // 6 *******
        8'b01111100, // 7   *****
        8'b01111000, // 8    ****
        8'b01110000, // 9     ***
        8'b01100000, // a      **
        8'b01000000, // b       *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x12
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00111100, // 3   ****
        8'b01111110, // 4  ******
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b01111110, // 8  ******
        8'b00111100, // 9   ****
        8'b00011000, // a    **
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x13
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100110, // 2  **  **
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b01100110, // 6  **  **
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b00000000, // 9
        8'b01100110, // a  **  **
        8'b01100110, // b  **  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x14
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2  *******
        8'b11011011, // 3 ** ** **
        8'b11011011, // 4 ** ** **
        8'b11011011, // 5 ** ** **
        8'b11011110, // 6  **** **
        8'b11011000, // 7    ** **
        8'b11011000, // 8    ** **
        8'b11011000, // 9    ** **
        8'b11011000, // a    ** **
        8'b11011000, // b    ** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x15
        8'b00000000, // 0
        8'b00111110, // 1  *****
        8'b01100011, // 2 **   **
        8'b00000110, // 3  **
        8'b00011100, // 4   ***
        8'b00110110, // 5  ** **
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b00110110, // 8  ** **
        8'b00011100, // 9   ***
        8'b00110000, // a     **
        8'b01100011, // b **   **
        8'b00111110, // c  *****
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x16
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b01111111, // 8 *******
        8'b01111111, // 9 *******
        8'b01111111, // a *******
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x17
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00111100, // 3   ****
        8'b01111110, // 4  ******
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b01111110, // 8  ******
        8'b00111100, // 9   ****
        8'b00011000, // a    **
        8'b01111110, // b  ******
        8'b00001100, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x18
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00111100, // 3   ****
        8'b01111110, // 4  ******
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x19
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b01111110, // 9  ******
        8'b00111100, // a   ****
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00011000, // 5    **
        8'b00110000, // 6     **
        8'b01111111, // 7 *******
        8'b00110000, // 8     **
        8'b00011000, // 9    **
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00001100, // 5   **
        8'b00000110, // 6  **
        8'b01111111, // 7 *******
        8'b00000110, // 8  **
        8'b00001100, // 9   **
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000011, // 6 **
        8'b00000011, // 7 **
        8'b00000011, // 8 **
        8'b01111111, // 9 *******
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00100100, // 5   *  *
        8'b01100110, // 6  **  **
        8'b11111111, // 7 ********
        8'b01100110, // 8  **  **
        8'b00100100, // 9   *  *
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00001000, // 4    *
        8'b00011100, // 5   ***
        8'b00011100, // 6   ***
        8'b00111110, // 7  *****
        8'b00111110, // 8  *****
        8'b01111111, // 9 *******
        8'b01111111, // a *******
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x1f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b01111111, // 4 *******
        8'b01111111, // 5 *******
        8'b00111110, // 6  *****
        8'b00111110, // 7  *****
        8'b00011100, // 8   ***
        8'b00011100, // 9   ***
        8'b00001000, // a    *
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x20
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x21
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00111100, // 3   ****
        8'b00111100, // 4   ****
        8'b00111100, // 5   ****
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00000000, // 9
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x22
        8'b00000000, // 0
        8'b01100110, // 1  **  **
        8'b01100110, // 2  **  **
        8'b01100110, // 3  **  **
        8'b00100100, // 4   *  *
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x23
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00110110, // 3  ** **
        8'b00110110, // 4  ** **
        8'b01111111, // 5 *******
        8'b00110110, // 6  ** **
        8'b00110110, // 7  ** **
        8'b00110110, // 8  ** **
        8'b01111111, // 9 *******
        8'b00110110, // a  ** **
        8'b00110110, // b  ** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x24
        8'b00011000, // 0     **
        8'b00011000, // 1     **
        8'b00111110, // 2   *****
        8'b01100011, // 3  **   **
        8'b01000011, // 4  **    *
        8'b00000011, // 5  **
        8'b00111110, // 6   *****
        8'b01100000, // 7       **
        8'b01100000, // 8       **
        8'b01100001, // 9  *    **
        8'b01100011, // a  **   **
        8'b00111110, // b   *****
        8'b00011000, // c     **
        8'b00011000, // d     **
        8'b00000000, // e
        8'b00000000, // f
         // code x25
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b01000011, // 4 **    *
        8'b01100011, // 5 **   **
        8'b00110000, // 6     **
        8'b00011000, // 7    **
        8'b00001100, // 8   **
        8'b00000110, // 9  **
        8'b01100011, // a **   **
        8'b01100001, // b *    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x26
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011100, // 2   ***
        8'b00110110, // 3  ** **
        8'b00110110, // 4  ** **
        8'b00011100, // 5   ***
        8'b01101110, // 6  *** **
        8'b00111011, // 7 ** ***
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b01101110, // b  *** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x27
        8'b00000000, // 0
        8'b00001100, // 1   **
        8'b00001100, // 2   **
        8'b00001100, // 3   **
        8'b00000110, // 4  **
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x28
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00110000, // 2     **
        8'b00011000, // 3    **
        8'b00001100, // 4   **
        8'b00001100, // 5   **
        8'b00001100, // 6   **
        8'b00001100, // 7   **
        8'b00001100, // 8   **
        8'b00001100, // 9   **
        8'b00011000, // a    **
        8'b00110000, // b     **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x29
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001100, // 2   **
        8'b00011000, // 3    **
        8'b00110000, // 4     **
        8'b00110000, // 5     **
        8'b00110000, // 6     **
        8'b00110000, // 7     **
        8'b00110000, // 8     **
        8'b00110000, // 9     **
        8'b00011000, // a    **
        8'b00001100, // b   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01100110, // 5  **  **
        8'b00111100, // 6   ****
        8'b11111111, // 7 ********
        8'b00111100, // 8   ****
        8'b01100110, // 9  **  **
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b01111110, // 7  ******
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00001100, // c   **
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b01111110, // 7  ******
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x2f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b01000000, // 4       *
        8'b01100000, // 5      **
        8'b00110000, // 6     **
        8'b00011000, // 7    **
        8'b00001100, // 8   **
        8'b00000110, // 9  **
        8'b00000011, // a **
        8'b00000001, // b *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x30
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01110011, // 5 **  ***
        8'b01111011, // 6 ** ****
        8'b01101111, // 7 **** **
        8'b01100111, // 8 ***  **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x31
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2
        8'b00011100, // 3
        8'b00011110, // 4    **
        8'b00011000, // 5   ***
        8'b00011000, // 6  ****
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b01111110, // b    **
        8'b00000000, // c    **
        8'b00000000, // d  ******
        8'b00000000, // e
        8'b00000000, // f
         // code x32
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100000, // 4      **
        8'b00110000, // 5     **
        8'b00011000, // 6    **
        8'b00001100, // 7   **
        8'b00000110, // 8  **
        8'b00000011, // 9 **
        8'b01100011, // a **   **
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x33
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100000, // 4      **
        8'b01100000, // 5      **
        8'b00111100, // 6   ****
        8'b01100000, // 7      **
        8'b01100000, // 8      **
        8'b01100000, // 9      **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x34
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00110000, // 2     **
        8'b00111000, // 3    ***
        8'b00111100, // 4   ****
        8'b00110110, // 5  ** **
        8'b00110011, // 6 **  **
        8'b01111111, // 7 *******
        8'b00110000, // 8     **
        8'b00110000, // 9     **
        8'b00110000, // a     **
        8'b01111000, // b    ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x35
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b00000011, // 3 **
        8'b00000011, // 4 **
        8'b00000011, // 5 **
        8'b00111111, // 6 ******
        8'b01100000, // 7      **
        8'b01100000, // 8      **
        8'b01100000, // 9      **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x36
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011100, // 2   ***
        8'b00000110, // 3  **
        8'b00000011, // 4 **
        8'b00000011, // 5 **
        8'b00111111, // 6 ******
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x37
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b01100011, // 3 **   **
        8'b01100000, // 4      **
        8'b01100000, // 5      **
        8'b00110000, // 6     **
        8'b00011000, // 7    **
        8'b00001100, // 8   **
        8'b00001100, // 9   **
        8'b00001100, // a   **
        8'b00001100, // b   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x38
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b00111110, // 6  *****
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x39
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111110, // 6  ******
        8'b01100000, // 7      **
        8'b01100000, // 8      **
        8'b01100000, // 9      **
        8'b00110000, // a     **
        8'b00011110, // b  ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00001100, // b   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b01100000, // 3      **
        8'b00110000, // 4     **
        8'b00011000, // 5    **
        8'b00001100, // 6   **
        8'b00000110, // 7  **
        8'b00001100, // 8   **
        8'b00011000, // 9    **
        8'b00110000, // a     **
        8'b01100000, // b      **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01111110, // 5  ******
        8'b00000000, // 6
        8'b00000000, // 7
        8'b01111110, // 8  ******
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000110, // 3  **
        8'b00001100, // 4   **
        8'b00011000, // 5    **
        8'b00110000, // 6     **
        8'b01100000, // 7      **
        8'b00110000, // 8     **
        8'b00011000, // 9    **
        8'b00001100, // a   **
        8'b00000110, // b  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x3f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b00110000, // 5     **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00000000, // 9
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x40
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111011, // 6 ** ****
        8'b01111011, // 7 ** ****
        8'b01111011, // 8 ** ****
        8'b00111011, // 9 ** ***
        8'b00000011, // a **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x41
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001000, // 2    *
        8'b00011100, // 3   ***
        8'b00110110, // 4  ** **
        8'b01100011, // 5 **   **
        8'b01100011, // 6 **   **
        8'b01111111, // 7 *******
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01100011, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x42
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111111, // 2 ******
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b00111110, // 6  *****
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b00111111, // b ******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x43
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b01100110, // 3  **  **
        8'b01000011, // 4 **    *
        8'b00000011, // 5 **
        8'b00000011, // 6 **
        8'b00000011, // 7 **
        8'b00000011, // 8 **
        8'b01000011, // 9 **    *
        8'b01100110, // a  **  **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x44
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011111, // 2 *****
        8'b00110110, // 3  ** **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b01100110, // 6  **  **
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b00110110, // a  ** **
        8'b00011111, // b *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x45
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b01100110, // 3  **  **
        8'b01000110, // 4  **   *
        8'b00010110, // 5  ** *
        8'b00011110, // 6  ****
        8'b00010110, // 7  ** *
        8'b00000110, // 8  **
        8'b01000110, // 9  **   *
        8'b01100110, // a  **  **
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x46
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b01100110, // 3  **  **
        8'b01000110, // 4  **   *
        8'b00010110, // 5  ** *
        8'b00011110, // 6  ****
        8'b00010110, // 7  ** *
        8'b00000110, // 8  **
        8'b00000110, // 9  **
        8'b00000110, // a  **
        8'b00001111, // b ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x47
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b01100110, // 3  **  **
        8'b01000011, // 4 **    *
        8'b00000011, // 5 **
        8'b00000011, // 6 **
        8'b01111011, // 7 ** ****
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100110, // a  **  **
        8'b01011100, // b   *** *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x48
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100011, // 2 **   **
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111111, // 6 *******
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01100011, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x49
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111000, // 2    ****
        8'b00110000, // 3     **
        8'b00110000, // 4     **
        8'b00110000, // 5     **
        8'b00110000, // 6     **
        8'b00110000, // 7     **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b00011110, // b  ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100111, // 2 ***  **
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b00110110, // 5  ** **
        8'b00011110, // 6  ****
        8'b00011110, // 7  ****
        8'b00110110, // 8  ** **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b01100111, // b ***  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001111, // 2 ****
        8'b00000110, // 3  **
        8'b00000110, // 4  **
        8'b00000110, // 5  **
        8'b00000110, // 6  **
        8'b00000110, // 7  **
        8'b00000110, // 8  **
        8'b01000110, // 9  **   *
        8'b01100110, // a  **  **
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000011, // 2 **    **
        8'b11100111, // 3 ***  ***
        8'b11111111, // 4 ********
        8'b11111111, // 5 ********
        8'b11011011, // 6 ** ** **
        8'b11000011, // 7 **    **
        8'b11000011, // 8 **    **
        8'b11000011, // 9 **    **
        8'b11000011, // a **    **
        8'b11000011, // b **    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100011, // 2 **   **
        8'b01100111, // 3 ***  **
        8'b01101111, // 4 **** **
        8'b01111111, // 5 *******
        8'b01111011, // 6 ** ****
        8'b01110011, // 7 **  ***
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01100011, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x4f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x50
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111111, // 2 ******
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b00111110, // 6  *****
        8'b00000110, // 7  **
        8'b00000110, // 8  **
        8'b00000110, // 9  **
        8'b00000110, // a  **
        8'b00001111, // b ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x510
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01101011, // 9 ** * **
        8'b01111011, // a ** ****
        8'b00111110, // b  *****
        8'b00110000, // c     **
        8'b01110000, // d     ***
        8'b00000000, // e
        8'b00000000, // f
         // code x52
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111111, // 2 ******
        8'b01100110, // 3  **  **
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b00111110, // 6  *****
        8'b00110110, // 7  ** **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b01100111, // b ***  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x53
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111110, // 2  *****
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b00000110, // 5  **
        8'b00011100, // 6   ***
        8'b00110000, // 7     **
        8'b01100000, // 8      **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x54
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111111, // 2 ********
        8'b11011011, // 3 ** ** **
        8'b10011001, // 4 *  **  *
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x55
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100011, // 2 **   **
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x56
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000011, // 2 **    **
        8'b11000011, // 3 **    **
        8'b11000011, // 4 **    **
        8'b11000011, // 5 **    **
        8'b11000011, // 6 **    **
        8'b11000011, // 7 **    **
        8'b11000011, // 8 **    **
        8'b01100110, // 9  **  **
        8'b00111100, // a   ****
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x57
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000011, // 2 **    **
        8'b11000011, // 3 **    **
        8'b11000011, // 4 **    **
        8'b11000011, // 5 **    **
        8'b11000011, // 6 **    **
        8'b11011011, // 7 ** ** **
        8'b11011011, // 8 ** ** **
        8'b11111111, // 9 ********
        8'b01100110, // a  **  **
        8'b01100110, // b  **  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
        
         // code x58
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000011, // 2 **    **
        8'b11000011, // 3 **    **
        8'b01100110, // 4  **  **
        8'b00111100, // 5   ****
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00111100, // 8   ****
        8'b01100110, // 9  **  **
        8'b11000011, // a **    **
        8'b11000011, // b **    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x59
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11000011, // 2 **    **
        8'b11000011, // 3 **    **
        8'b11000011, // 4 **    **
        8'b01100110, // 5  **  **
        8'b00111100, // 6   ****
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111111, // 2 ********
        8'b11000011, // 3 **    **
        8'b01100001, // 4 *    **
        8'b00110000, // 5     **
        8'b00011000, // 6    **
        8'b00001100, // 7   **
        8'b00000110, // 8  **
        8'b10000011, // 9 **     *
        8'b11000011, // a **    **
        8'b11111111, // b ********
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b00001100, // 3   **
        8'b00001100, // 4   **
        8'b00001100, // 5   **
        8'b00001100, // 6   **
        8'b00001100, // 7   **
        8'b00001100, // 8   **
        8'b00001100, // 9   **
        8'b00001100, // a   **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000001, // 3 *
        8'b00000011, // 4 **
        8'b00000111, // 5 ***
        8'b00001110, // 6  ***
        8'b00011100, // 7   ***
        8'b00111000, // 8    ***
        8'b01110000, // 9     ***
        8'b01100000, // a      **
        8'b01000000, // b       *
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b00110000, // 3     **
        8'b00110000, // 4     **
        8'b00110000, // 5     **
        8'b00110000, // 6     **
        8'b00110000, // 7     **
        8'b00110000, // 8     **
        8'b00110000, // 9     **
        8'b00110000, // a     **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5e
        8'b00001000, // 0    *
        8'b00011100, // 1   ***
        8'b00110110, // 2  ** **
        8'b01100011, // 3 **   **
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x5f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b11111111, // d ********
        8'b00000000, // e
        8'b00000000, // f
         // code x60
        8'b00001100, // 0   **
        8'b00001100, // 1   **
        8'b00011000, // 2    **
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x61
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00011110, // 5  ****
        8'b00110000, // 6     **
        8'b00111110, // 7  *****
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b01101110, // b  *** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x62
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000111, // 2  ***
        8'b00000110, // 3   **
        8'b00000110, // 4   **
        8'b00011110, // 5   ****
        8'b00110110, // 6   ** **
        8'b01100110, // 7   **  **
        8'b01100110, // 8   **  **
        8'b01100110, // 9   **  **
        8'b01100110, // a   **  **
        8'b00111110, // b   *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x63
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111110, // 5  *****
        8'b01100011, // 6 **   **
        8'b00000011, // 7 **
        8'b00000011, // 8 **
        8'b00000011, // 9 **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x64
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111000, // 2    ***
        8'b00110000, // 3     **
        8'b00110000, // 4     **
        8'b00111100, // 5   ****
        8'b00110110, // 6  ** **
        8'b00110011, // 7 **  **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b01101110, // b  *** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x65
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111110, // 5  *****
        8'b01100011, // 6 **   **
        8'b01111111, // 7 *******
        8'b00000011, // 8 **
        8'b00000011, // 9 **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x66
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011100, // 2   ***
        8'b00110110, // 3  ** **
        8'b00100110, // 4  **  *
        8'b00000110, // 5  **
        8'b00001111, // 6 ****
        8'b00000110, // 7  **
        8'b00000110, // 8  **
        8'b00000110, // 9  **
        8'b00000110, // a  **
        8'b00001111, // b ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x67
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01101110, // 5  *** **
        8'b00110011, // 6 **  **
        8'b00110011, // 7 **  **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b00111110, // b  *****
        8'b00110000, // c     **
        8'b00110011, // d **  **
        8'b00011110, // e  ****
        8'b00000000, // f
         // code x68
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000111, // 2 ***
        8'b00000110, // 3  **
        8'b00000110, // 4  **
        8'b00110110, // 5  ** **
        8'b01101110, // 6  *** **
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b01100111, // b ***  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x69
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00011000, // 3    **
        8'b00000000, // 4
        8'b00011100, // 5   ***
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x6a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100000, // 2      **
        8'b01100000, // 3      **
        8'b00000000, // 4
        8'b01110000, // 5     ***
        8'b01100000, // 6      **
        8'b01100000, // 7      **
        8'b01100000, // 8      **
        8'b01100000, // 9      **
        8'b01100000, // a      **
        8'b01100000, // b      **
        8'b01100110, // c  **  **
        8'b01100110, // d  **  **
        8'b00111100, // e   ****
        8'b00000000, // f
         // code x6b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000111, // 2 ***
        8'b00000110, // 3  **
        8'b00000110, // 4  **
        8'b01100110, // 5  **  **
        8'b00110110, // 6  ** **
        8'b00011110, // 7  ****
        8'b00011110, // 8  ****
        8'b00110110, // 9  ** **
        8'b01100110, // a  **  **
        8'b01100111, // b ***  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x6c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011100, // 2   ***
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00111100, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x6d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01100111, // 5 ***  **
        8'b11111111, // 6 ********
        8'b11011011, // 7 ** ** **
        8'b11011011, // 8 ** ** **
        8'b11011011, // 9 ** ** **
        8'b11011011, // a ** ** **
        8'b11011011, // b ** ** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x6e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111011, // 5 ** ***
        8'b01100110, // 6  **  **
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b01100110, // b  **  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x6f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111110, // 5  *****
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x70
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111011, // 5 ** ***
        8'b01100110, // 6  **  **
        8'b01100110, // 7  **  **
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b00111110, // b  *****
        8'b00000110, // c  **
        8'b00000110, // d  **
        8'b00001111, // e ****
        8'b00000000, // f
         // code x71
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01101110, // 5  *** **
        8'b00110011, // 6 **  **
        8'b00110011, // 7 **  **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b00111110, // b  *****
        8'b00110000, // c     **
        8'b00110000, // d     **
        8'b01111000, // e    ****
        8'b00000000, // f
         // code x72
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111011, // 5 ** ***
        8'b01101110, // 6  *** **
        8'b01100110, // 7  **  **
        8'b00000110, // 8  **
        8'b00000110, // 9  **
        8'b00000110, // a  **
        8'b00001111, // b ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x73
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00111110, // 5  *****
        8'b01100011, // 6 **   **
        8'b00000110, // 7  **
        8'b00011100, // 8   ***
        8'b00110000, // 9     **
        8'b01100011, // a **   **
        8'b00111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x74
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001000, // 2    *
        8'b00001100, // 3   **
        8'b00001100, // 4   **
        8'b00111111, // 5 ******
        8'b00001100, // 6   **
        8'b00001100, // 7   **
        8'b00001100, // 8   **
        8'b00001100, // 9   **
        8'b01101100, // a   ** **
        8'b00111000, // b    ***
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x75
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b00110011, // 5 **  **
        8'b00110011, // 6 **  **
        8'b00110011, // 7 **  **
        8'b00110011, // 8 **  **
        8'b00110011, // 9 **  **
        8'b00110011, // a **  **
        8'b01101110, // b  *** **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x76
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b11000011, // 5 **    **
        8'b11000011, // 6 **    **
        8'b11000011, // 7 **    **
        8'b11000011, // 8 **    **
        8'b01100110, // 9  **  **
        8'b00111100, // a   ****
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x77
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b11000011, // 5 **    **
        8'b11000011, // 6 **    **
        8'b11000011, // 7 **    **
        8'b11011011, // 8 ** ** **
        8'b11011011, // 9 ** ** **
        8'b11111111, // a ********
        8'b01100110, // b  **  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x78
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b11000011, // 5 **    **
        8'b01100110, // 6  **  **
        8'b00111100, // 7   ****
        8'b00011000, // 8    **
        8'b00111100, // 9   ****
        8'b01100110, // a  **  **
        8'b11000011, // b **    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x79
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01100011, // 5 **   **
        8'b01100011, // 6 **   **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01111110, // b  ******
        8'b01100000, // c      **
        8'b00110000, // d     **
        8'b00011111, // e *****
        8'b00000000, // f
         // code x7a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00000000, // 4
        8'b01111111, // 5 *******
        8'b00110011, // 6 **  **
        8'b00011000, // 7    **
        8'b00001100, // 8   **
        8'b00000110, // 9  **
        8'b01100011, // a **   **
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x7b
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01110000, // 2     ***
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00001110, // 6  ***
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b01110000, // b     ***
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x7c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00011000, // 2    **
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00000000, // 6
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x7d
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00001110, // 2  ***
        8'b00011000, // 3    **
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b01110000, // 6     ***
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00001110, // b  ***
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x7e
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01101110, // 2  *** **
        8'b00111011, // 3 ** ***
        8'b00000000, // 4
        8'b00000000, // 5
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00000000, // 9
        8'b00000000, // a
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
         // code x7f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00001000, // 4    *
        8'b00011100, // 5   ***
        8'b00110110, // 6  ** **
        8'b01100011, // 7 **   **
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01111111, // a *******
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000  // f
        };

	assign data = ROM[addr];

endmodule  